magic
tech sky130A
magscale 1 2
timestamp 1672326805
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1640 178848 117552
<< metal2 >>
rect 2962 0 3018 800
rect 8574 0 8630 800
rect 14186 0 14242 800
rect 19798 0 19854 800
rect 25410 0 25466 800
rect 31022 0 31078 800
rect 36634 0 36690 800
rect 42246 0 42302 800
rect 47858 0 47914 800
rect 53470 0 53526 800
rect 59082 0 59138 800
rect 64694 0 64750 800
rect 70306 0 70362 800
rect 75918 0 75974 800
rect 81530 0 81586 800
rect 87142 0 87198 800
rect 92754 0 92810 800
rect 98366 0 98422 800
rect 103978 0 104034 800
rect 109590 0 109646 800
rect 115202 0 115258 800
rect 120814 0 120870 800
rect 126426 0 126482 800
rect 132038 0 132094 800
rect 137650 0 137706 800
rect 143262 0 143318 800
rect 148874 0 148930 800
rect 154486 0 154542 800
rect 160098 0 160154 800
rect 165710 0 165766 800
rect 171322 0 171378 800
rect 176934 0 176990 800
<< obsm2 >>
rect 2964 856 176988 117541
rect 3074 734 8518 856
rect 8686 734 14130 856
rect 14298 734 19742 856
rect 19910 734 25354 856
rect 25522 734 30966 856
rect 31134 734 36578 856
rect 36746 734 42190 856
rect 42358 734 47802 856
rect 47970 734 53414 856
rect 53582 734 59026 856
rect 59194 734 64638 856
rect 64806 734 70250 856
rect 70418 734 75862 856
rect 76030 734 81474 856
rect 81642 734 87086 856
rect 87254 734 92698 856
rect 92866 734 98310 856
rect 98478 734 103922 856
rect 104090 734 109534 856
rect 109702 734 115146 856
rect 115314 734 120758 856
rect 120926 734 126370 856
rect 126538 734 131982 856
rect 132150 734 137594 856
rect 137762 734 143206 856
rect 143374 734 148818 856
rect 148986 734 154430 856
rect 154598 734 160042 856
rect 160210 734 165654 856
rect 165822 734 171266 856
rect 171434 734 176878 856
<< obsm3 >>
rect 4210 2075 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 43299 7379 43365 13293
<< labels >>
rlabel metal2 s 47858 0 47914 800 6 clk
port 1 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 clken
port 2 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 in[0]
port 3 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 in[1]
port 4 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 in[2]
port 5 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 in[3]
port 6 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 in[4]
port 7 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 in[5]
port 8 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 in[6]
port 9 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 in[7]
port 10 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 ld
port 11 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 ld1
port 12 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 ld2
port 13 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 ld3
port 14 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 ld4
port 15 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 out[0]
port 16 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 out[10]
port 17 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 out[11]
port 18 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 out[12]
port 19 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 out[13]
port 20 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 out[14]
port 21 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 out[15]
port 22 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 out[1]
port 23 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 out[2]
port 24 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 out[3]
port 25 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 out[4]
port 26 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 out[5]
port 27 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 out[6]
port 28 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 out[7]
port 29 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 out[8]
port 30 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 out[9]
port 31 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 rst
port 32 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9350412
string GDS_FILE /home/sky/MPW8/IIT_Indore_MAC_MPW8/openlane/mac/runs/22_12_29_06_57/results/signoff/mac.magic.gds
string GDS_START 500640
<< end >>

