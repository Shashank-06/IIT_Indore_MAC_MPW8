// This is the unpowered netlist.
module mac (clk,
    clken,
    ld,
    ld1,
    ld2,
    ld3,
    ld4,
    rst,
    in,
    io_oeb,
    out);
 input clk;
 input clken;
 input ld;
 input ld1;
 input ld2;
 input ld3;
 input ld4;
 input rst;
 input [7:0] in;
 output [15:0] io_oeb;
 output [15:0] out;

 wire \A1.x[0] ;
 wire \A1.x[1] ;
 wire \A1.x[2] ;
 wire \A1.x[3] ;
 wire \A1.x[4] ;
 wire \A1.x[5] ;
 wire \A1.x[6] ;
 wire \A1.x[7] ;
 wire \I1.out[0] ;
 wire \I1.out[1] ;
 wire \I1.out[2] ;
 wire \I1.out[3] ;
 wire \I1.out[4] ;
 wire \I1.out[5] ;
 wire \I1.out[6] ;
 wire \I1.out[7] ;
 wire \I2.out[0] ;
 wire \I2.out[1] ;
 wire \I2.out[2] ;
 wire \I2.out[3] ;
 wire \I2.out[4] ;
 wire \I2.out[5] ;
 wire \I2.out[6] ;
 wire \I2.out[7] ;
 wire \I3.out[0] ;
 wire \I3.out[1] ;
 wire \I3.out[2] ;
 wire \I3.out[3] ;
 wire \I3.out[4] ;
 wire \I3.out[5] ;
 wire \I3.out[6] ;
 wire \I3.out[7] ;
 wire \I4.out[0] ;
 wire \I4.out[1] ;
 wire \I4.out[2] ;
 wire \I4.out[3] ;
 wire \I4.out[4] ;
 wire \I4.out[5] ;
 wire \I4.out[6] ;
 wire \I4.out[7] ;
 wire \P1.in[0] ;
 wire \P1.in[10] ;
 wire \P1.in[11] ;
 wire \P1.in[12] ;
 wire \P1.in[13] ;
 wire \P1.in[14] ;
 wire \P1.in[15] ;
 wire \P1.in[1] ;
 wire \P1.in[2] ;
 wire \P1.in[3] ;
 wire \P1.in[4] ;
 wire \P1.in[5] ;
 wire \P1.in[6] ;
 wire \P1.in[7] ;
 wire \P1.in[8] ;
 wire \P1.in[9] ;
 wire \P1.qq[10] ;
 wire \P1.qq[11] ;
 wire \P1.qq[12] ;
 wire \P1.qq[13] ;
 wire \P1.qq[14] ;
 wire \P1.qq[15] ;
 wire \P1.qq[8] ;
 wire \P1.qq[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire net26;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire \m1.a[0] ;
 wire \m1.a[1] ;
 wire \m1.a[2] ;
 wire \m1.a[3] ;
 wire \m1.a[4] ;
 wire \m1.a[5] ;
 wire \m1.a[6] ;
 wire \m1.a[7] ;
 wire \m1.b[0] ;
 wire \m1.b[1] ;
 wire \m1.b[2] ;
 wire \m1.b[3] ;
 wire \m1.b[4] ;
 wire \m1.b[5] ;
 wire \m1.b[6] ;
 wire \m1.b[7] ;
 wire \m1.multa_reg[0] ;
 wire \m1.multa_reg[10] ;
 wire \m1.multa_reg[11] ;
 wire \m1.multa_reg[12] ;
 wire \m1.multa_reg[13] ;
 wire \m1.multa_reg[14] ;
 wire \m1.multa_reg[15] ;
 wire \m1.multa_reg[1] ;
 wire \m1.multa_reg[2] ;
 wire \m1.multa_reg[3] ;
 wire \m1.multa_reg[4] ;
 wire \m1.multa_reg[5] ;
 wire \m1.multa_reg[6] ;
 wire \m1.multa_reg[7] ;
 wire \m1.multa_reg[8] ;
 wire \m1.multa_reg[9] ;
 wire \m1.out[0] ;
 wire \m1.out[10] ;
 wire \m1.out[11] ;
 wire \m1.out[12] ;
 wire \m1.out[13] ;
 wire \m1.out[14] ;
 wire \m1.out[15] ;
 wire \m1.out[16] ;
 wire \m1.out[1] ;
 wire \m1.out[2] ;
 wire \m1.out[3] ;
 wire \m1.out[4] ;
 wire \m1.out[5] ;
 wire \m1.out[6] ;
 wire \m1.out[7] ;
 wire \m1.out[8] ;
 wire \m1.out[9] ;
 wire \m2.a[0] ;
 wire \m2.a[1] ;
 wire \m2.a[2] ;
 wire \m2.a[3] ;
 wire \m2.a[4] ;
 wire \m2.a[5] ;
 wire \m2.a[6] ;
 wire \m2.a[7] ;
 wire \m2.b[0] ;
 wire \m2.b[1] ;
 wire \m2.b[2] ;
 wire \m2.b[3] ;
 wire \m2.b[4] ;
 wire \m2.b[5] ;
 wire \m2.b[6] ;
 wire \m2.b[7] ;
 wire \m2.multa_reg[0] ;
 wire \m2.multa_reg[10] ;
 wire \m2.multa_reg[11] ;
 wire \m2.multa_reg[12] ;
 wire \m2.multa_reg[13] ;
 wire \m2.multa_reg[14] ;
 wire \m2.multa_reg[15] ;
 wire \m2.multa_reg[1] ;
 wire \m2.multa_reg[2] ;
 wire \m2.multa_reg[3] ;
 wire \m2.multa_reg[4] ;
 wire \m2.multa_reg[5] ;
 wire \m2.multa_reg[6] ;
 wire \m2.multa_reg[7] ;
 wire \m2.multa_reg[8] ;
 wire \m2.multa_reg[9] ;
 wire \m2.out[0] ;
 wire \m2.out[10] ;
 wire \m2.out[11] ;
 wire \m2.out[12] ;
 wire \m2.out[13] ;
 wire \m2.out[14] ;
 wire \m2.out[15] ;
 wire \m2.out[16] ;
 wire \m2.out[1] ;
 wire \m2.out[2] ;
 wire \m2.out[3] ;
 wire \m2.out[4] ;
 wire \m2.out[5] ;
 wire \m2.out[6] ;
 wire \m2.out[7] ;
 wire \m2.out[8] ;
 wire \m2.out[9] ;
 wire net42;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net48;

 sky130_fd_sc_hd__buf_2 _1239_ (.A(\m2.a[7] ),
    .X(_0696_));
 sky130_fd_sc_hd__buf_2 _1240_ (.A(\m2.a[6] ),
    .X(_0697_));
 sky130_fd_sc_hd__buf_2 _1241_ (.A(\m2.b[7] ),
    .X(_0698_));
 sky130_fd_sc_hd__buf_2 _1242_ (.A(\m2.b[6] ),
    .X(_0699_));
 sky130_fd_sc_hd__nand4_1 _1243_ (.A(_0696_),
    .B(_0697_),
    .C(_0698_),
    .D(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__a22o_1 _1244_ (.A1(_0697_),
    .A2(_0698_),
    .B1(_0699_),
    .B2(_0696_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_2 _1245_ (.A(\m2.b[5] ),
    .X(_0702_));
 sky130_fd_sc_hd__buf_2 _1246_ (.A(\m2.a[5] ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(_0703_),
    .B(_0698_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand2_1 _1248_ (.A(_0697_),
    .B(_0699_),
    .Y(_0705_));
 sky130_fd_sc_hd__buf_2 _1249_ (.A(\m2.b[4] ),
    .X(_0706_));
 sky130_fd_sc_hd__and2_1 _1250_ (.A(_0697_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__and3_1 _1251_ (.A(_0696_),
    .B(_0702_),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(_0705_),
    .A1(_0699_),
    .S(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__xor2_1 _1253_ (.A(_0704_),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__and3_1 _1254_ (.A(_0696_),
    .B(_0702_),
    .C(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__and3_1 _1255_ (.A(_0700_),
    .B(_0701_),
    .C(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0700_),
    .A2(_0701_),
    .B1(_0711_),
    .Y(_0713_));
 sky130_fd_sc_hd__or2_1 _1257_ (.A(_0712_),
    .B(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__o2bb2ai_1 _1258_ (.A1_N(_0699_),
    .A2_N(_0708_),
    .B1(_0709_),
    .B2(_0704_),
    .Y(_0715_));
 sky130_fd_sc_hd__and2b_1 _1259_ (.A_N(_0714_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__and3_1 _1260_ (.A(_0696_),
    .B(_0698_),
    .C(_0705_),
    .X(_0717_));
 sky130_fd_sc_hd__o21a_1 _1261_ (.A1(_0712_),
    .A2(_0716_),
    .B1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__a21oi_1 _1262_ (.A1(_0696_),
    .A2(_0702_),
    .B1(_0710_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_1 _1263_ (.A(_0711_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__a22oi_1 _1264_ (.A1(_0697_),
    .A2(_0702_),
    .B1(_0706_),
    .B2(_0696_),
    .Y(_0721_));
 sky130_fd_sc_hd__or2_1 _1265_ (.A(_0708_),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_4 _1266_ (.A(\m2.b[3] ),
    .X(_0723_));
 sky130_fd_sc_hd__a21o_1 _1267_ (.A1(_0696_),
    .A2(_0723_),
    .B1(_0707_),
    .X(_0724_));
 sky130_fd_sc_hd__and3_1 _1268_ (.A(\m2.a[7] ),
    .B(_0723_),
    .C(_0707_),
    .X(_0725_));
 sky130_fd_sc_hd__a31o_1 _1269_ (.A1(_0703_),
    .A2(_0702_),
    .A3(_0724_),
    .B1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__a21oi_1 _1270_ (.A1(_0703_),
    .A2(_0699_),
    .B1(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__and3_1 _1271_ (.A(_0703_),
    .B(_0699_),
    .C(_0726_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1272_ (.A(_0727_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__buf_2 _1273_ (.A(\m2.a[4] ),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(_0730_),
    .B(_0698_),
    .Y(_0731_));
 sky130_fd_sc_hd__xnor2_1 _1275_ (.A(_0729_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__and2b_1 _1276_ (.A_N(_0722_),
    .B(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__and2_1 _1277_ (.A(_0720_),
    .B(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__a31oi_2 _1278_ (.A1(_0730_),
    .A2(_0698_),
    .A3(_0729_),
    .B1(_0728_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _1279_ (.A(_0720_),
    .B(_0733_),
    .Y(_0736_));
 sky130_fd_sc_hd__nor2_1 _1280_ (.A(_0734_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__and2b_1 _1281_ (.A_N(_0735_),
    .B(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__xnor2_1 _1282_ (.A(_0715_),
    .B(_0714_),
    .Y(_0739_));
 sky130_fd_sc_hd__o21a_1 _1283_ (.A1(_0734_),
    .A2(_0738_),
    .B1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__inv_2 _1284_ (.A(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _1285_ (.A(_0730_),
    .B(_0702_),
    .Y(_0742_));
 sky130_fd_sc_hd__a22oi_1 _1286_ (.A1(_0703_),
    .A2(_0706_),
    .B1(_0723_),
    .B2(_0697_),
    .Y(_0743_));
 sky130_fd_sc_hd__and3_1 _1287_ (.A(_0703_),
    .B(_0723_),
    .C(_0707_),
    .X(_0744_));
 sky130_fd_sc_hd__o21bai_1 _1288_ (.A1(_0742_),
    .A2(_0743_),
    .B1_N(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__and3_1 _1289_ (.A(_0730_),
    .B(_0699_),
    .C(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__clkbuf_4 _1290_ (.A(\m2.a[3] ),
    .X(_0747_));
 sky130_fd_sc_hd__a21oi_1 _1291_ (.A1(_0730_),
    .A2(_0699_),
    .B1(_0745_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _1292_ (.A(_0748_),
    .B(_0746_),
    .Y(_0749_));
 sky130_fd_sc_hd__and3_1 _1293_ (.A(_0747_),
    .B(_0698_),
    .C(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__or2_1 _1294_ (.A(_0746_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__buf_2 _1295_ (.A(\m2.b[2] ),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _1296_ (.A(\m2.b[1] ),
    .X(_0753_));
 sky130_fd_sc_hd__and4_1 _1297_ (.A(\m2.a[7] ),
    .B(_0697_),
    .C(_0752_),
    .D(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _1298_ (.A(_0743_),
    .B(_0744_),
    .Y(_0755_));
 sky130_fd_sc_hd__xnor2_1 _1299_ (.A(_0742_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_1 _1300_ (.A(_0697_),
    .B(_0753_),
    .Y(_0757_));
 sky130_fd_sc_hd__and3_1 _1301_ (.A(_0696_),
    .B(_0752_),
    .C(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__and2_1 _1302_ (.A(_0756_),
    .B(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _1303_ (.A(_0703_),
    .B(_0702_),
    .Y(_0760_));
 sky130_fd_sc_hd__and2b_1 _1304_ (.A_N(_0725_),
    .B(_0724_),
    .X(_0761_));
 sky130_fd_sc_hd__xnor2_1 _1305_ (.A(_0760_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__o21a_1 _1306_ (.A1(_0754_),
    .A2(_0759_),
    .B1(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__a21oi_1 _1307_ (.A1(_0747_),
    .A2(_0698_),
    .B1(_0749_),
    .Y(_0764_));
 sky130_fd_sc_hd__nor3_1 _1308_ (.A(_0754_),
    .B(_0759_),
    .C(_0762_),
    .Y(_0765_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(_0763_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__nor3_1 _1310_ (.A(_0764_),
    .B(_0750_),
    .C(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(_0722_),
    .B(_0732_),
    .Y(_0768_));
 sky130_fd_sc_hd__o21a_1 _1312_ (.A1(_0763_),
    .A2(_0767_),
    .B1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__nor3_1 _1313_ (.A(_0763_),
    .B(_0767_),
    .C(_0768_),
    .Y(_0770_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a21o_1 _1315_ (.A1(_0751_),
    .A2(_0771_),
    .B1(_0769_),
    .X(_0772_));
 sky130_fd_sc_hd__xnor2_1 _1316_ (.A(_0735_),
    .B(_0737_),
    .Y(_0773_));
 sky130_fd_sc_hd__and2_1 _1317_ (.A(_0772_),
    .B(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0747_),
    .B(\m2.b[5] ),
    .Y(_0775_));
 sky130_fd_sc_hd__a22oi_1 _1319_ (.A1(_0730_),
    .A2(_0706_),
    .B1(_0723_),
    .B2(_0703_),
    .Y(_0776_));
 sky130_fd_sc_hd__and4_1 _1320_ (.A(_0703_),
    .B(_0730_),
    .C(_0706_),
    .D(\m2.b[3] ),
    .X(_0777_));
 sky130_fd_sc_hd__o21bai_1 _1321_ (.A1(_0775_),
    .A2(_0776_),
    .B1_N(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__and2_1 _1322_ (.A(_0747_),
    .B(\m2.b[6] ),
    .X(_0779_));
 sky130_fd_sc_hd__nor2_1 _1323_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__and2_1 _1324_ (.A(_0778_),
    .B(_0779_),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__buf_2 _1326_ (.A(\m2.a[2] ),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _1327_ (.A(_0783_),
    .B(\m2.b[7] ),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1328_ (.A(_0782_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__and2_1 _1329_ (.A(_0782_),
    .B(_0784_),
    .X(_0786_));
 sky130_fd_sc_hd__or2_1 _1330_ (.A(_0785_),
    .B(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _1331_ (.A(\m2.a[5] ),
    .B(_0752_),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _1332_ (.A1(\m2.a[6] ),
    .A2(\m2.b[1] ),
    .B1(\m2.b[0] ),
    .B2(\m2.a[7] ),
    .X(_0789_));
 sky130_fd_sc_hd__buf_2 _1333_ (.A(\m2.b[0] ),
    .X(_0790_));
 sky130_fd_sc_hd__nand4_1 _1334_ (.A(\m2.a[7] ),
    .B(\m2.a[6] ),
    .C(_0753_),
    .D(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__a21bo_1 _1335_ (.A1(_0788_),
    .A2(_0789_),
    .B1_N(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__a22oi_1 _1336_ (.A1(_0697_),
    .A2(_0752_),
    .B1(_0753_),
    .B2(\m2.a[7] ),
    .Y(_0793_));
 sky130_fd_sc_hd__nor2_1 _1337_ (.A(_0754_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__nor2_1 _1338_ (.A(_0776_),
    .B(_0777_),
    .Y(_0795_));
 sky130_fd_sc_hd__xnor2_1 _1339_ (.A(_0775_),
    .B(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__xor2_1 _1340_ (.A(_0792_),
    .B(_0794_),
    .X(_0797_));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0796_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__a21bo_1 _1342_ (.A1(_0792_),
    .A2(_0794_),
    .B1_N(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__xnor2_1 _1343_ (.A(_0756_),
    .B(_0758_),
    .Y(_0800_));
 sky130_fd_sc_hd__xor2_1 _1344_ (.A(_0799_),
    .B(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__or2b_1 _1345_ (.A(_0800_),
    .B_N(_0799_),
    .X(_0802_));
 sky130_fd_sc_hd__o21a_1 _1346_ (.A1(_0787_),
    .A2(_0801_),
    .B1(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _1347_ (.A(_0764_),
    .B(_0750_),
    .Y(_0804_));
 sky130_fd_sc_hd__xnor2_1 _1348_ (.A(_0804_),
    .B(_0766_),
    .Y(_0805_));
 sky130_fd_sc_hd__or2b_1 _1349_ (.A(_0803_),
    .B_N(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__xnor2_1 _1350_ (.A(_0803_),
    .B(_0805_),
    .Y(_0807_));
 sky130_fd_sc_hd__o21ai_1 _1351_ (.A1(_0781_),
    .A2(_0786_),
    .B1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__xnor2_1 _1352_ (.A(_0751_),
    .B(_0771_),
    .Y(_0809_));
 sky130_fd_sc_hd__a21oi_1 _1353_ (.A1(_0806_),
    .A2(_0808_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__or3_1 _1354_ (.A(_0781_),
    .B(_0786_),
    .C(_0807_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_0808_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__buf_2 _1356_ (.A(\m2.a[1] ),
    .X(_0813_));
 sky130_fd_sc_hd__a22oi_1 _1357_ (.A1(_0747_),
    .A2(_0706_),
    .B1(\m2.b[3] ),
    .B2(_0730_),
    .Y(_0814_));
 sky130_fd_sc_hd__and4_1 _1358_ (.A(_0730_),
    .B(_0747_),
    .C(\m2.b[4] ),
    .D(\m2.b[3] ),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(_0814_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__a31o_1 _1360_ (.A1(_0783_),
    .A2(_0702_),
    .A3(_0816_),
    .B1(_0815_),
    .X(_0817_));
 sky130_fd_sc_hd__a21oi_1 _1361_ (.A1(_0783_),
    .A2(\m2.b[6] ),
    .B1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__and3_1 _1362_ (.A(_0783_),
    .B(\m2.b[6] ),
    .C(_0817_),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_1 _1363_ (.A(_0818_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a31o_1 _1364_ (.A1(_0813_),
    .A2(_0698_),
    .A3(_0820_),
    .B1(_0819_),
    .X(_0821_));
 sky130_fd_sc_hd__nand3_1 _1365_ (.A(_0791_),
    .B(_0788_),
    .C(_0789_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_1 _1366_ (.A(\m2.a[4] ),
    .B(_0752_),
    .Y(_0823_));
 sky130_fd_sc_hd__a22oi_2 _1367_ (.A1(\m2.a[5] ),
    .A2(\m2.b[1] ),
    .B1(\m2.b[0] ),
    .B2(\m2.a[6] ),
    .Y(_0824_));
 sky130_fd_sc_hd__and4_1 _1368_ (.A(\m2.a[6] ),
    .B(\m2.a[5] ),
    .C(\m2.b[1] ),
    .D(\m2.b[0] ),
    .X(_0825_));
 sky130_fd_sc_hd__o21bai_1 _1369_ (.A1(_0823_),
    .A2(_0824_),
    .B1_N(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a21o_1 _1370_ (.A1(_0791_),
    .A2(_0789_),
    .B1(_0788_),
    .X(_0827_));
 sky130_fd_sc_hd__nand3_1 _1371_ (.A(_0822_),
    .B(_0826_),
    .C(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _1372_ (.A(_0783_),
    .B(_0702_),
    .Y(_0829_));
 sky130_fd_sc_hd__xnor2_1 _1373_ (.A(_0829_),
    .B(_0816_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21o_1 _1374_ (.A1(_0822_),
    .A2(_0827_),
    .B1(_0826_),
    .X(_0831_));
 sky130_fd_sc_hd__nand3_1 _1375_ (.A(_0828_),
    .B(_0830_),
    .C(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0828_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__or2_1 _1377_ (.A(_0796_),
    .B(_0797_),
    .X(_0834_));
 sky130_fd_sc_hd__and3_1 _1378_ (.A(_0798_),
    .B(_0833_),
    .C(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0813_),
    .B(\m2.b[7] ),
    .Y(_0836_));
 sky130_fd_sc_hd__xor2_1 _1380_ (.A(_0820_),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nand2_1 _1381_ (.A(_0798_),
    .B(_0834_),
    .Y(_0838_));
 sky130_fd_sc_hd__xnor2_1 _1382_ (.A(_0833_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__and2b_1 _1383_ (.A_N(_0837_),
    .B(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__xor2_1 _1384_ (.A(_0787_),
    .B(_0801_),
    .X(_0841_));
 sky130_fd_sc_hd__or3_1 _1385_ (.A(_0835_),
    .B(_0840_),
    .C(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__o21ai_1 _1386_ (.A1(_0835_),
    .A2(_0840_),
    .B1(_0841_),
    .Y(_0843_));
 sky130_fd_sc_hd__a21bo_1 _1387_ (.A1(_0821_),
    .A2(_0842_),
    .B1_N(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__or2b_1 _1388_ (.A(_0812_),
    .B_N(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(_0843_),
    .B(_0842_),
    .X(_0846_));
 sky130_fd_sc_hd__xnor2_1 _1390_ (.A(_0821_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_0813_),
    .B(\m2.b[5] ),
    .Y(_0848_));
 sky130_fd_sc_hd__a22oi_1 _1392_ (.A1(\m2.a[2] ),
    .A2(_0706_),
    .B1(\m2.b[3] ),
    .B2(_0747_),
    .Y(_0849_));
 sky130_fd_sc_hd__and4_1 _1393_ (.A(\m2.a[3] ),
    .B(\m2.a[2] ),
    .C(\m2.b[4] ),
    .D(\m2.b[3] ),
    .X(_0850_));
 sky130_fd_sc_hd__nor2_1 _1394_ (.A(_0849_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__xnor2_1 _1395_ (.A(_0848_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__or3_1 _1396_ (.A(_0825_),
    .B(_0823_),
    .C(_0824_),
    .X(_0853_));
 sky130_fd_sc_hd__o21ai_1 _1397_ (.A1(_0825_),
    .A2(_0824_),
    .B1(_0823_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _1398_ (.A(\m2.a[3] ),
    .B(\m2.b[2] ),
    .Y(_0855_));
 sky130_fd_sc_hd__a22oi_2 _1399_ (.A1(\m2.a[4] ),
    .A2(\m2.b[1] ),
    .B1(\m2.b[0] ),
    .B2(\m2.a[5] ),
    .Y(_0856_));
 sky130_fd_sc_hd__and4_1 _1400_ (.A(\m2.a[5] ),
    .B(\m2.a[4] ),
    .C(\m2.b[1] ),
    .D(\m2.b[0] ),
    .X(_0857_));
 sky130_fd_sc_hd__o21bai_1 _1401_ (.A1(_0855_),
    .A2(_0856_),
    .B1_N(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a21o_1 _1402_ (.A1(_0853_),
    .A2(_0854_),
    .B1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__nand3_1 _1403_ (.A(_0853_),
    .B(_0858_),
    .C(_0854_),
    .Y(_0860_));
 sky130_fd_sc_hd__a21bo_1 _1404_ (.A1(_0852_),
    .A2(_0859_),
    .B1_N(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__a21o_1 _1405_ (.A1(_0828_),
    .A2(_0831_),
    .B1(_0830_),
    .X(_0862_));
 sky130_fd_sc_hd__nand3_1 _1406_ (.A(_0832_),
    .B(_0861_),
    .C(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__o21bai_1 _1407_ (.A1(_0848_),
    .A2(_0849_),
    .B1_N(_0850_),
    .Y(_0864_));
 sky130_fd_sc_hd__and2_1 _1408_ (.A(_0813_),
    .B(\m2.b[6] ),
    .X(_0865_));
 sky130_fd_sc_hd__nor2_1 _1409_ (.A(_0864_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__and2_1 _1410_ (.A(_0864_),
    .B(_0865_),
    .X(_0867_));
 sky130_fd_sc_hd__nor2_1 _1411_ (.A(_0866_),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__buf_2 _1412_ (.A(\m2.a[0] ),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _1413_ (.A(_0869_),
    .B(\m2.b[7] ),
    .Y(_0870_));
 sky130_fd_sc_hd__xnor2_1 _1414_ (.A(_0868_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21o_1 _1415_ (.A1(_0832_),
    .A2(_0862_),
    .B1(_0861_),
    .X(_0872_));
 sky130_fd_sc_hd__nand3_1 _1416_ (.A(_0863_),
    .B(_0871_),
    .C(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__and2_1 _1417_ (.A(_0863_),
    .B(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__xor2_1 _1418_ (.A(_0837_),
    .B(_0839_),
    .X(_0875_));
 sky130_fd_sc_hd__o21ba_1 _1419_ (.A1(_0866_),
    .A2(_0870_),
    .B1_N(_0867_),
    .X(_0876_));
 sky130_fd_sc_hd__xor2_1 _1420_ (.A(_0874_),
    .B(_0875_),
    .X(_0877_));
 sky130_fd_sc_hd__or2b_1 _1421_ (.A(_0876_),
    .B_N(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__o21ai_1 _1422_ (.A1(_0874_),
    .A2(_0875_),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__or2b_1 _1423_ (.A(_0847_),
    .B_N(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__nand3_1 _1424_ (.A(_0860_),
    .B(_0852_),
    .C(_0859_),
    .Y(_0881_));
 sky130_fd_sc_hd__a22o_1 _1425_ (.A1(\m2.a[1] ),
    .A2(\m2.b[4] ),
    .B1(\m2.b[3] ),
    .B2(\m2.a[2] ),
    .X(_0882_));
 sky130_fd_sc_hd__nand4_1 _1426_ (.A(\m2.a[2] ),
    .B(\m2.a[1] ),
    .C(\m2.b[4] ),
    .D(\m2.b[3] ),
    .Y(_0883_));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(\m2.a[0] ),
    .B(\m2.b[5] ),
    .X(_0884_));
 sky130_fd_sc_hd__a21oi_1 _1428_ (.A1(_0882_),
    .A2(_0883_),
    .B1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__and3_1 _1429_ (.A(_0884_),
    .B(_0882_),
    .C(_0883_),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _1430_ (.A(_0885_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__or3_1 _1431_ (.A(_0857_),
    .B(_0855_),
    .C(_0856_),
    .X(_0888_));
 sky130_fd_sc_hd__o21ai_1 _1432_ (.A1(_0857_),
    .A2(_0856_),
    .B1(_0855_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_1 _1433_ (.A(\m2.a[2] ),
    .B(_0752_),
    .Y(_0890_));
 sky130_fd_sc_hd__a22oi_2 _1434_ (.A1(_0747_),
    .A2(\m2.b[1] ),
    .B1(_0790_),
    .B2(\m2.a[4] ),
    .Y(_0891_));
 sky130_fd_sc_hd__and4_1 _1435_ (.A(\m2.a[4] ),
    .B(\m2.a[3] ),
    .C(\m2.b[1] ),
    .D(\m2.b[0] ),
    .X(_0892_));
 sky130_fd_sc_hd__o21bai_1 _1436_ (.A1(_0890_),
    .A2(_0891_),
    .B1_N(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__a21o_1 _1437_ (.A1(_0888_),
    .A2(_0889_),
    .B1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nand3_1 _1438_ (.A(_0888_),
    .B(_0893_),
    .C(_0889_),
    .Y(_0895_));
 sky130_fd_sc_hd__a21bo_1 _1439_ (.A1(_0887_),
    .A2(_0894_),
    .B1_N(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__a21o_1 _1440_ (.A1(_0860_),
    .A2(_0859_),
    .B1(_0852_),
    .X(_0897_));
 sky130_fd_sc_hd__and3_1 _1441_ (.A(_0881_),
    .B(_0896_),
    .C(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__and4_1 _1442_ (.A(_0783_),
    .B(_0813_),
    .C(_0706_),
    .D(_0723_),
    .X(_0899_));
 sky130_fd_sc_hd__o211a_1 _1443_ (.A1(_0899_),
    .A2(_0886_),
    .B1(_0869_),
    .C1(\m2.b[6] ),
    .X(_0900_));
 sky130_fd_sc_hd__a211oi_1 _1444_ (.A1(_0869_),
    .A2(\m2.b[6] ),
    .B1(_0899_),
    .C1(_0886_),
    .Y(_0901_));
 sky130_fd_sc_hd__or2_1 _1445_ (.A(_0900_),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a21oi_1 _1446_ (.A1(_0881_),
    .A2(_0897_),
    .B1(_0896_),
    .Y(_0903_));
 sky130_fd_sc_hd__nor3_1 _1447_ (.A(_0898_),
    .B(_0902_),
    .C(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a21o_1 _1448_ (.A1(_0863_),
    .A2(_0872_),
    .B1(_0871_),
    .X(_0905_));
 sky130_fd_sc_hd__o211a_1 _1449_ (.A1(_0898_),
    .A2(_0904_),
    .B1(_0905_),
    .C1(_0873_),
    .X(_0906_));
 sky130_fd_sc_hd__a211oi_1 _1450_ (.A1(_0873_),
    .A2(_0905_),
    .B1(_0904_),
    .C1(_0898_),
    .Y(_0907_));
 sky130_fd_sc_hd__or3b_1 _1451_ (.A(_0906_),
    .B(_0907_),
    .C_N(_0900_),
    .X(_0908_));
 sky130_fd_sc_hd__or2b_1 _1452_ (.A(_0906_),
    .B_N(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__xnor2_1 _1453_ (.A(_0876_),
    .B(_0877_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _1454_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand3_1 _1455_ (.A(_0895_),
    .B(_0887_),
    .C(_0894_),
    .Y(_0912_));
 sky130_fd_sc_hd__a22o_1 _1456_ (.A1(\m2.a[0] ),
    .A2(_0706_),
    .B1(_0723_),
    .B2(_0813_),
    .X(_0913_));
 sky130_fd_sc_hd__and4_1 _1457_ (.A(\m2.a[1] ),
    .B(\m2.a[0] ),
    .C(\m2.b[4] ),
    .D(\m2.b[3] ),
    .X(_0914_));
 sky130_fd_sc_hd__inv_2 _1458_ (.A(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(_0913_),
    .B(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__or3_1 _1460_ (.A(_0892_),
    .B(_0890_),
    .C(_0891_),
    .X(_0917_));
 sky130_fd_sc_hd__o21ai_1 _1461_ (.A1(_0892_),
    .A2(_0891_),
    .B1(_0890_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _1462_ (.A(_0813_),
    .B(_0752_),
    .Y(_0919_));
 sky130_fd_sc_hd__a22oi_1 _1463_ (.A1(_0783_),
    .A2(_0753_),
    .B1(_0790_),
    .B2(_0747_),
    .Y(_0920_));
 sky130_fd_sc_hd__and4_1 _1464_ (.A(\m2.a[3] ),
    .B(\m2.a[2] ),
    .C(\m2.b[1] ),
    .D(_0790_),
    .X(_0921_));
 sky130_fd_sc_hd__o21bai_1 _1465_ (.A1(_0919_),
    .A2(_0920_),
    .B1_N(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__a21o_1 _1466_ (.A1(_0917_),
    .A2(_0918_),
    .B1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__and3_1 _1467_ (.A(_0917_),
    .B(_0922_),
    .C(_0918_),
    .X(_0924_));
 sky130_fd_sc_hd__a21o_1 _1468_ (.A1(_0916_),
    .A2(_0923_),
    .B1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(_0895_),
    .A2(_0894_),
    .B1(_0887_),
    .X(_0926_));
 sky130_fd_sc_hd__and3_1 _1470_ (.A(_0912_),
    .B(_0925_),
    .C(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__a21oi_1 _1471_ (.A1(_0912_),
    .A2(_0926_),
    .B1(_0925_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor3_1 _1472_ (.A(_0915_),
    .B(_0927_),
    .C(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__o21ai_1 _1473_ (.A1(_0898_),
    .A2(_0903_),
    .B1(_0902_),
    .Y(_0930_));
 sky130_fd_sc_hd__or3_1 _1474_ (.A(_0898_),
    .B(_0902_),
    .C(_0903_),
    .X(_0931_));
 sky130_fd_sc_hd__o211a_1 _1475_ (.A1(_0927_),
    .A2(_0929_),
    .B1(_0930_),
    .C1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__o21bai_1 _1476_ (.A1(_0906_),
    .A2(_0907_),
    .B1_N(_0900_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand3_1 _1477_ (.A(_0908_),
    .B(_0932_),
    .C(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__and3_1 _1478_ (.A(_0908_),
    .B(_0932_),
    .C(_0933_),
    .X(_0935_));
 sky130_fd_sc_hd__a21oi_1 _1479_ (.A1(_0908_),
    .A2(_0933_),
    .B1(_0932_),
    .Y(_0936_));
 sky130_fd_sc_hd__a211oi_1 _1480_ (.A1(_0931_),
    .A2(_0930_),
    .B1(_0929_),
    .C1(_0927_),
    .Y(_0937_));
 sky130_fd_sc_hd__and4_1 _1481_ (.A(_0783_),
    .B(\m2.a[1] ),
    .C(_0753_),
    .D(_0790_),
    .X(_0938_));
 sky130_fd_sc_hd__a22oi_1 _1482_ (.A1(\m2.a[1] ),
    .A2(_0753_),
    .B1(_0790_),
    .B2(_0783_),
    .Y(_0939_));
 sky130_fd_sc_hd__and4bb_1 _1483_ (.A_N(_0938_),
    .B_N(_0939_),
    .C(\m2.a[0] ),
    .D(_0752_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(_0938_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_0921_),
    .B(_0920_),
    .Y(_0942_));
 sky130_fd_sc_hd__xnor2_1 _1486_ (.A(_0919_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__and2b_1 _1487_ (.A_N(_0941_),
    .B(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__xnor2_1 _1488_ (.A(_0941_),
    .B(_0943_),
    .Y(_0945_));
 sky130_fd_sc_hd__and3_1 _1489_ (.A(_0869_),
    .B(_0723_),
    .C(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__and2b_1 _1490_ (.A_N(_0924_),
    .B(_0923_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _1491_ (.A(_0916_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__o21ai_2 _1492_ (.A1(_0944_),
    .A2(_0946_),
    .B1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__o21a_1 _1493_ (.A1(_0927_),
    .A2(_0928_),
    .B1(_0915_),
    .X(_0950_));
 sky130_fd_sc_hd__or2_1 _1494_ (.A(_0929_),
    .B(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__o22a_1 _1495_ (.A1(_0932_),
    .A2(_0937_),
    .B1(_0949_),
    .B2(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__and4_1 _1496_ (.A(_0813_),
    .B(_0869_),
    .C(_0753_),
    .D(_0790_),
    .X(_0953_));
 sky130_fd_sc_hd__o2bb2a_1 _1497_ (.A1_N(_0869_),
    .A2_N(_0752_),
    .B1(_0938_),
    .B2(_0939_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2_1 _1498_ (.A(_0940_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__and2_1 _1499_ (.A(_0953_),
    .B(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__nand2_1 _1500_ (.A(_0869_),
    .B(_0723_),
    .Y(_0957_));
 sky130_fd_sc_hd__xnor2_1 _1501_ (.A(_0957_),
    .B(_0945_),
    .Y(_0958_));
 sky130_fd_sc_hd__and2_1 _1502_ (.A(_0956_),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__or3_1 _1503_ (.A(_0948_),
    .B(_0944_),
    .C(_0946_),
    .X(_0960_));
 sky130_fd_sc_hd__nand3_1 _1504_ (.A(_0949_),
    .B(_0959_),
    .C(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__or2_1 _1505_ (.A(_0951_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__or4_1 _1506_ (.A(_0932_),
    .B(_0937_),
    .C(_0949_),
    .D(_0951_),
    .X(_0963_));
 sky130_fd_sc_hd__o21ai_1 _1507_ (.A1(_0952_),
    .A2(_0962_),
    .B1(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__or3b_1 _1508_ (.A(_0935_),
    .B(_0936_),
    .C_N(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__xnor2_1 _1509_ (.A(_0909_),
    .B(_0910_),
    .Y(_0966_));
 sky130_fd_sc_hd__a21o_1 _1510_ (.A1(_0934_),
    .A2(_0965_),
    .B1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__xor2_1 _1511_ (.A(_0879_),
    .B(_0847_),
    .X(_0968_));
 sky130_fd_sc_hd__a21o_1 _1512_ (.A1(_0911_),
    .A2(_0967_),
    .B1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__xor2_1 _1513_ (.A(_0844_),
    .B(_0812_),
    .X(_0970_));
 sky130_fd_sc_hd__a21o_1 _1514_ (.A1(_0880_),
    .A2(_0969_),
    .B1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__and3_1 _1515_ (.A(_0806_),
    .B(_0808_),
    .C(_0809_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_1 _1516_ (.A(_0810_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__a21oi_1 _1517_ (.A1(_0845_),
    .A2(_0971_),
    .B1(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__or2_1 _1518_ (.A(_0772_),
    .B(_0773_),
    .X(_0975_));
 sky130_fd_sc_hd__and2b_1 _1519_ (.A_N(_0774_),
    .B(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__o21a_1 _1520_ (.A1(_0810_),
    .A2(_0974_),
    .B1(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__or3_1 _1521_ (.A(_0734_),
    .B(_0738_),
    .C(_0739_),
    .X(_0978_));
 sky130_fd_sc_hd__and2_1 _1522_ (.A(_0741_),
    .B(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__o21ai_1 _1523_ (.A1(_0774_),
    .A2(_0977_),
    .B1(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__or3_1 _1524_ (.A(_0712_),
    .B(_0716_),
    .C(_0717_),
    .X(_0981_));
 sky130_fd_sc_hd__and2b_1 _1525_ (.A_N(_0718_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a21boi_1 _1526_ (.A1(_0741_),
    .A2(_0980_),
    .B1_N(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__buf_4 _1527_ (.A(net1),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_4 _1528_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(_0985_),
    .B(_0700_),
    .Y(_0986_));
 sky130_fd_sc_hd__o32a_1 _1530_ (.A1(_0718_),
    .A2(_0983_),
    .A3(_0986_),
    .B1(_0985_),
    .B2(\m2.multa_reg[15] ),
    .X(_0259_));
 sky130_fd_sc_hd__inv_2 _1531_ (.A(net1),
    .Y(_0987_));
 sky130_fd_sc_hd__clkbuf_4 _1532_ (.A(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__and3b_1 _1533_ (.A_N(_0982_),
    .B(_0741_),
    .C(_0980_),
    .X(_0989_));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_0988_),
    .B(\m2.multa_reg[14] ),
    .Y(_0990_));
 sky130_fd_sc_hd__o31ai_1 _1535_ (.A1(_0988_),
    .A2(_0983_),
    .A3(_0989_),
    .B1(_0990_),
    .Y(_0258_));
 sky130_fd_sc_hd__clkbuf_4 _1536_ (.A(_0987_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_4 _1537_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_4 _1538_ (.A(_0984_),
    .X(_0993_));
 sky130_fd_sc_hd__or3_1 _1539_ (.A(_0979_),
    .B(_0774_),
    .C(_0977_),
    .X(_0994_));
 sky130_fd_sc_hd__and3_1 _1540_ (.A(_0993_),
    .B(_0980_),
    .C(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a21o_1 _1541_ (.A1(_0992_),
    .A2(\m2.multa_reg[13] ),
    .B1(_0995_),
    .X(_0257_));
 sky130_fd_sc_hd__nor3_1 _1542_ (.A(_0976_),
    .B(_0810_),
    .C(_0974_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_0977_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\m2.multa_reg[12] ),
    .A1(_0997_),
    .S(_0993_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0998_),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _1546_ (.A(_0973_),
    .B(_0845_),
    .C(_0971_),
    .X(_0999_));
 sky130_fd_sc_hd__or3_1 _1547_ (.A(_0987_),
    .B(_0974_),
    .C(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__a21bo_1 _1548_ (.A1(_0992_),
    .A2(\m2.multa_reg[11] ),
    .B1_N(_1000_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _1549_ (.A(_0970_),
    .B(_0880_),
    .C(_0969_),
    .X(_1001_));
 sky130_fd_sc_hd__or3b_1 _1550_ (.A(_1001_),
    .B(_0987_),
    .C_N(_0971_),
    .X(_1002_));
 sky130_fd_sc_hd__a21bo_1 _1551_ (.A1(_0992_),
    .A2(\m2.multa_reg[10] ),
    .B1_N(_1002_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _1552_ (.A(_0968_),
    .B(_0911_),
    .C(_0967_),
    .X(_1003_));
 sky130_fd_sc_hd__or3b_1 _1553_ (.A(_1003_),
    .B(_0987_),
    .C_N(_0969_),
    .X(_1004_));
 sky130_fd_sc_hd__a21bo_1 _1554_ (.A1(_0992_),
    .A2(\m2.multa_reg[9] ),
    .B1_N(_1004_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _1555_ (.A(_0966_),
    .B(_0934_),
    .C(_0965_),
    .X(_1005_));
 sky130_fd_sc_hd__or3b_1 _1556_ (.A(_1005_),
    .B(_0987_),
    .C_N(_0967_),
    .X(_1006_));
 sky130_fd_sc_hd__a21bo_1 _1557_ (.A1(_0992_),
    .A2(\m2.multa_reg[8] ),
    .B1_N(_1006_),
    .X(_0252_));
 sky130_fd_sc_hd__o21bai_1 _1558_ (.A1(_0935_),
    .A2(_0936_),
    .B1_N(_0964_),
    .Y(_1007_));
 sky130_fd_sc_hd__and2_1 _1559_ (.A(_0991_),
    .B(\m2.multa_reg[7] ),
    .X(_1008_));
 sky130_fd_sc_hd__a31o_1 _1560_ (.A1(_0985_),
    .A2(_0965_),
    .A3(_1007_),
    .B1(_1008_),
    .X(_0251_));
 sky130_fd_sc_hd__nor4_1 _1561_ (.A(_0932_),
    .B(_0937_),
    .C(_0949_),
    .D(_0951_),
    .Y(_1009_));
 sky130_fd_sc_hd__nor2_1 _1562_ (.A(_1009_),
    .B(_0952_),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_1 _1563_ (.A(_1010_),
    .B(_0962_),
    .Y(_1011_));
 sky130_fd_sc_hd__buf_4 _1564_ (.A(net1),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(\m2.multa_reg[6] ),
    .A1(_1011_),
    .S(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _1566_ (.A(_1013_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _1567_ (.A(_0949_),
    .B(_0961_),
    .Y(_1014_));
 sky130_fd_sc_hd__xnor2_1 _1568_ (.A(_0951_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(\m2.multa_reg[5] ),
    .A1(_1015_),
    .S(_1012_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _1570_ (.A(_1016_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _1571_ (.A1(_0949_),
    .A2(_0960_),
    .B1(_0959_),
    .X(_1017_));
 sky130_fd_sc_hd__and3_1 _1572_ (.A(_0993_),
    .B(_0961_),
    .C(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__a21o_1 _1573_ (.A1(_0992_),
    .A2(\m2.multa_reg[4] ),
    .B1(_1018_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _1574_ (.A(_0956_),
    .B(_0958_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _1575_ (.A(_0959_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(\m2.multa_reg[3] ),
    .A1(_1020_),
    .S(_1012_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _1577_ (.A(_1021_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _1578_ (.A(_0953_),
    .B(_0955_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _1579_ (.A(_0991_),
    .B(_0956_),
    .Y(_1023_));
 sky130_fd_sc_hd__a22o_1 _1580_ (.A1(_0988_),
    .A2(\m2.multa_reg[2] ),
    .B1(_1022_),
    .B2(_1023_),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _1581_ (.A1(_0869_),
    .A2(_0753_),
    .B1(_0790_),
    .B2(_0813_),
    .X(_1024_));
 sky130_fd_sc_hd__nor2_1 _1582_ (.A(_0991_),
    .B(_0953_),
    .Y(_1025_));
 sky130_fd_sc_hd__a22o_1 _1583_ (.A1(_0988_),
    .A2(\m2.multa_reg[1] ),
    .B1(_1024_),
    .B2(_1025_),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _1584_ (.A(_0993_),
    .B(_0869_),
    .C(_0790_),
    .X(_1026_));
 sky130_fd_sc_hd__a21o_1 _1585_ (.A1(_0992_),
    .A2(\m2.multa_reg[0] ),
    .B1(_1026_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_2 _1586_ (.A(\m1.a[7] ),
    .X(_1027_));
 sky130_fd_sc_hd__buf_2 _1587_ (.A(\m1.a[6] ),
    .X(_1028_));
 sky130_fd_sc_hd__buf_2 _1588_ (.A(\m1.b[7] ),
    .X(_1029_));
 sky130_fd_sc_hd__buf_2 _1589_ (.A(\m1.b[6] ),
    .X(_1030_));
 sky130_fd_sc_hd__and4_1 _1590_ (.A(_1027_),
    .B(_1028_),
    .C(_1029_),
    .D(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__a22oi_1 _1591_ (.A1(_1028_),
    .A2(_1029_),
    .B1(_1030_),
    .B2(_1027_),
    .Y(_1032_));
 sky130_fd_sc_hd__nor2_1 _1592_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__buf_2 _1593_ (.A(\m1.b[5] ),
    .X(_1034_));
 sky130_fd_sc_hd__buf_2 _1594_ (.A(\m1.a[5] ),
    .X(_1035_));
 sky130_fd_sc_hd__nand2_1 _1595_ (.A(_1035_),
    .B(_1029_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand2_1 _1596_ (.A(_1028_),
    .B(_1030_),
    .Y(_1037_));
 sky130_fd_sc_hd__clkbuf_4 _1597_ (.A(\m1.b[4] ),
    .X(_1038_));
 sky130_fd_sc_hd__and2_1 _1598_ (.A(_1028_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nand3_1 _1599_ (.A(_1027_),
    .B(_1034_),
    .C(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__clkinv_2 _1600_ (.A(\m1.b[6] ),
    .Y(_1041_));
 sky130_fd_sc_hd__or2_1 _1601_ (.A(_1041_),
    .B(_1040_),
    .X(_1042_));
 sky130_fd_sc_hd__a21bo_1 _1602_ (.A1(_1037_),
    .A2(_1040_),
    .B1_N(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__and2_1 _1603_ (.A(_1036_),
    .B(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nor2_1 _1604_ (.A(_1036_),
    .B(_1043_),
    .Y(_1045_));
 sky130_fd_sc_hd__nor2_1 _1605_ (.A(_1044_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__and3_1 _1606_ (.A(_1027_),
    .B(_1034_),
    .C(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__inv_2 _1607_ (.A(_1045_),
    .Y(_1048_));
 sky130_fd_sc_hd__xnor2_1 _1608_ (.A(_1033_),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__a21oi_1 _1609_ (.A1(_1042_),
    .A2(_1048_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__a21o_1 _1610_ (.A1(_1033_),
    .A2(_1047_),
    .B1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__and3_1 _1611_ (.A(_1027_),
    .B(_1029_),
    .C(_1037_),
    .X(_1052_));
 sky130_fd_sc_hd__a21o_1 _1612_ (.A1(_1051_),
    .A2(_1052_),
    .B1(_1031_),
    .X(_1053_));
 sky130_fd_sc_hd__a21oi_1 _1613_ (.A1(_1027_),
    .A2(_1034_),
    .B1(_1046_),
    .Y(_1054_));
 sky130_fd_sc_hd__nor2_1 _1614_ (.A(_1047_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__a22o_1 _1615_ (.A1(_1028_),
    .A2(_1034_),
    .B1(_1038_),
    .B2(_1027_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_2 _1616_ (.A(\m1.a[4] ),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_4 _1617_ (.A(\m1.b[3] ),
    .X(_1058_));
 sky130_fd_sc_hd__a21o_1 _1618_ (.A1(_1027_),
    .A2(_1058_),
    .B1(_1039_),
    .X(_1059_));
 sky130_fd_sc_hd__and3_1 _1619_ (.A(\m1.a[7] ),
    .B(_1058_),
    .C(_1039_),
    .X(_1060_));
 sky130_fd_sc_hd__a31o_1 _1620_ (.A1(_1035_),
    .A2(_1034_),
    .A3(_1059_),
    .B1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__a21oi_1 _1621_ (.A1(_1035_),
    .A2(_1030_),
    .B1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__and3_1 _1622_ (.A(_1035_),
    .B(_1030_),
    .C(_1061_),
    .X(_1063_));
 sky130_fd_sc_hd__nor2_1 _1623_ (.A(_1062_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__a21oi_1 _1624_ (.A1(_1057_),
    .A2(_1029_),
    .B1(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__and3_1 _1625_ (.A(_1057_),
    .B(_1029_),
    .C(_1064_),
    .X(_1066_));
 sky130_fd_sc_hd__nor2_1 _1626_ (.A(_1065_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__and3_1 _1627_ (.A(_1040_),
    .B(_1056_),
    .C(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _1628_ (.A(_1055_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__or2_1 _1629_ (.A(_1055_),
    .B(_1068_),
    .X(_1070_));
 sky130_fd_sc_hd__and2_1 _1630_ (.A(_1069_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_1 _1631_ (.A1(_1063_),
    .A2(_1066_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__and3_1 _1632_ (.A(_1042_),
    .B(_1048_),
    .C(_1049_),
    .X(_1073_));
 sky130_fd_sc_hd__or2_1 _1633_ (.A(_1050_),
    .B(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__a21o_1 _1634_ (.A1(_1069_),
    .A2(_1072_),
    .B1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__buf_2 _1635_ (.A(\m1.b[2] ),
    .X(_1076_));
 sky130_fd_sc_hd__buf_2 _1636_ (.A(\m1.b[1] ),
    .X(_1077_));
 sky130_fd_sc_hd__and4_1 _1637_ (.A(\m1.a[7] ),
    .B(_1028_),
    .C(_1076_),
    .D(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _1638_ (.A(_1057_),
    .B(_1034_),
    .Y(_1079_));
 sky130_fd_sc_hd__a22oi_1 _1639_ (.A1(_1035_),
    .A2(_1038_),
    .B1(_1058_),
    .B2(_1028_),
    .Y(_1080_));
 sky130_fd_sc_hd__and3_1 _1640_ (.A(_1035_),
    .B(_1058_),
    .C(_1039_),
    .X(_1081_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__xnor2_1 _1642_ (.A(_1079_),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__nand2_1 _1643_ (.A(_1028_),
    .B(_1077_),
    .Y(_1084_));
 sky130_fd_sc_hd__and3_1 _1644_ (.A(_1027_),
    .B(_1076_),
    .C(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _1645_ (.A(_1083_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__nand2_1 _1646_ (.A(_1035_),
    .B(_1034_),
    .Y(_1087_));
 sky130_fd_sc_hd__and2b_1 _1647_ (.A_N(_1060_),
    .B(_1059_),
    .X(_1088_));
 sky130_fd_sc_hd__xnor2_1 _1648_ (.A(_1087_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__o21a_1 _1649_ (.A1(_1078_),
    .A2(_1086_),
    .B1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__buf_2 _1650_ (.A(\m1.a[3] ),
    .X(_1091_));
 sky130_fd_sc_hd__o21bai_1 _1651_ (.A1(_1079_),
    .A2(_1080_),
    .B1_N(_1081_),
    .Y(_1092_));
 sky130_fd_sc_hd__a21oi_1 _1652_ (.A1(_1057_),
    .A2(_1030_),
    .B1(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__and3_1 _1653_ (.A(_1057_),
    .B(_1030_),
    .C(_1092_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _1654_ (.A(_1093_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__a21oi_1 _1655_ (.A1(_1091_),
    .A2(_1029_),
    .B1(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__and3_1 _1656_ (.A(_1091_),
    .B(_1029_),
    .C(_1095_),
    .X(_1097_));
 sky130_fd_sc_hd__nor3_1 _1657_ (.A(_1078_),
    .B(_1086_),
    .C(_1089_),
    .Y(_1098_));
 sky130_fd_sc_hd__or2_1 _1658_ (.A(_1090_),
    .B(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__nor3_1 _1659_ (.A(_1096_),
    .B(_1097_),
    .C(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__a21oi_1 _1660_ (.A1(_1040_),
    .A2(_1056_),
    .B1(_1067_),
    .Y(_1101_));
 sky130_fd_sc_hd__nor2_1 _1661_ (.A(_1068_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__o21ai_1 _1662_ (.A1(_1090_),
    .A2(_1100_),
    .B1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__or2_1 _1663_ (.A(_1094_),
    .B(_1097_),
    .X(_1104_));
 sky130_fd_sc_hd__or3_1 _1664_ (.A(_1090_),
    .B(_1100_),
    .C(_1102_),
    .X(_1105_));
 sky130_fd_sc_hd__and2_1 _1665_ (.A(_1103_),
    .B(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_1 _1666_ (.A(_1104_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__or3_1 _1667_ (.A(_1063_),
    .B(_1066_),
    .C(_1071_),
    .X(_1108_));
 sky130_fd_sc_hd__nand2_1 _1668_ (.A(_1072_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a21o_1 _1669_ (.A1(_1103_),
    .A2(_1107_),
    .B1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__xnor2_2 _1670_ (.A(_1104_),
    .B(_1106_),
    .Y(_1111_));
 sky130_fd_sc_hd__a22oi_1 _1671_ (.A1(_1057_),
    .A2(_1038_),
    .B1(_1058_),
    .B2(_1035_),
    .Y(_1112_));
 sky130_fd_sc_hd__and4_1 _1672_ (.A(_1035_),
    .B(_1057_),
    .C(\m1.b[4] ),
    .D(\m1.b[3] ),
    .X(_1113_));
 sky130_fd_sc_hd__nor2_1 _1673_ (.A(_1112_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__a31o_1 _1674_ (.A1(_1091_),
    .A2(_1034_),
    .A3(_1114_),
    .B1(_1113_),
    .X(_1115_));
 sky130_fd_sc_hd__and2_1 _1675_ (.A(_1091_),
    .B(\m1.b[6] ),
    .X(_1116_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__buf_2 _1677_ (.A(\m1.a[2] ),
    .X(_1118_));
 sky130_fd_sc_hd__nand2_1 _1678_ (.A(_1118_),
    .B(\m1.b[7] ),
    .Y(_1119_));
 sky130_fd_sc_hd__and2_1 _1679_ (.A(_1115_),
    .B(_1116_),
    .X(_1120_));
 sky130_fd_sc_hd__o21bai_1 _1680_ (.A1(_1117_),
    .A2(_1119_),
    .B1_N(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__or2_1 _1681_ (.A(_1117_),
    .B(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__xnor2_1 _1682_ (.A(_1122_),
    .B(_1119_),
    .Y(_1123_));
 sky130_fd_sc_hd__and2_1 _1683_ (.A(\m1.a[5] ),
    .B(_1076_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_2 _1684_ (.A(\m1.b[0] ),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _1685_ (.A1(\m1.a[6] ),
    .A2(\m1.b[1] ),
    .B1(_1125_),
    .B2(\m1.a[7] ),
    .X(_1126_));
 sky130_fd_sc_hd__nand4_1 _1686_ (.A(\m1.a[7] ),
    .B(\m1.a[6] ),
    .C(_1077_),
    .D(_1125_),
    .Y(_1127_));
 sky130_fd_sc_hd__a21bo_1 _1687_ (.A1(_1124_),
    .A2(_1126_),
    .B1_N(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a22oi_1 _1688_ (.A1(_1028_),
    .A2(_1076_),
    .B1(_1077_),
    .B2(\m1.a[7] ),
    .Y(_1129_));
 sky130_fd_sc_hd__nor2_1 _1689_ (.A(_1078_),
    .B(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_1 _1690_ (.A(_1091_),
    .B(\m1.b[5] ),
    .Y(_1131_));
 sky130_fd_sc_hd__xnor2_1 _1691_ (.A(_1131_),
    .B(_1114_),
    .Y(_1132_));
 sky130_fd_sc_hd__xor2_1 _1692_ (.A(_1128_),
    .B(_1130_),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__a21bo_1 _1694_ (.A1(_1128_),
    .A2(_1130_),
    .B1_N(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__xnor2_1 _1695_ (.A(_1083_),
    .B(_1085_),
    .Y(_1136_));
 sky130_fd_sc_hd__xor2_1 _1696_ (.A(_1135_),
    .B(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__or2b_1 _1697_ (.A(_1136_),
    .B_N(_1135_),
    .X(_1138_));
 sky130_fd_sc_hd__o21a_1 _1698_ (.A1(_1123_),
    .A2(_1137_),
    .B1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_1 _1699_ (.A(_1096_),
    .B(_1097_),
    .Y(_1140_));
 sky130_fd_sc_hd__xnor2_1 _1700_ (.A(_1140_),
    .B(_1099_),
    .Y(_1141_));
 sky130_fd_sc_hd__xnor2_1 _1701_ (.A(_1139_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__or2b_1 _1702_ (.A(_1139_),
    .B_N(_1141_),
    .X(_1143_));
 sky130_fd_sc_hd__a21bo_1 _1703_ (.A1(_1121_),
    .A2(_1142_),
    .B1_N(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__or2b_1 _1704_ (.A(_1111_),
    .B_N(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__nand3_1 _1705_ (.A(_1127_),
    .B(_1124_),
    .C(_1126_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(\m1.a[4] ),
    .B(\m1.b[2] ),
    .Y(_1147_));
 sky130_fd_sc_hd__a22oi_2 _1707_ (.A1(\m1.a[5] ),
    .A2(\m1.b[1] ),
    .B1(\m1.b[0] ),
    .B2(\m1.a[6] ),
    .Y(_1148_));
 sky130_fd_sc_hd__and4_1 _1708_ (.A(\m1.a[6] ),
    .B(\m1.a[5] ),
    .C(\m1.b[1] ),
    .D(\m1.b[0] ),
    .X(_1149_));
 sky130_fd_sc_hd__o21bai_1 _1709_ (.A1(_1147_),
    .A2(_1148_),
    .B1_N(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__a21o_1 _1710_ (.A1(_1127_),
    .A2(_1126_),
    .B1(_1124_),
    .X(_1151_));
 sky130_fd_sc_hd__nand3_1 _1711_ (.A(_1146_),
    .B(_1150_),
    .C(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_1118_),
    .B(\m1.b[5] ),
    .Y(_1153_));
 sky130_fd_sc_hd__a22oi_1 _1713_ (.A1(_1091_),
    .A2(_1038_),
    .B1(\m1.b[3] ),
    .B2(_1057_),
    .Y(_1154_));
 sky130_fd_sc_hd__and4_1 _1714_ (.A(_1057_),
    .B(_1091_),
    .C(\m1.b[4] ),
    .D(\m1.b[3] ),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _1715_ (.A(_1154_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__xnor2_1 _1716_ (.A(_1153_),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__a21o_1 _1717_ (.A1(_1146_),
    .A2(_1151_),
    .B1(_1150_),
    .X(_1158_));
 sky130_fd_sc_hd__nand3_1 _1718_ (.A(_1152_),
    .B(_1157_),
    .C(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _1719_ (.A(_1152_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__or2_1 _1720_ (.A(_1132_),
    .B(_1133_),
    .X(_1161_));
 sky130_fd_sc_hd__and3_1 _1721_ (.A(_1134_),
    .B(_1160_),
    .C(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__a31o_1 _1722_ (.A1(_1118_),
    .A2(_1034_),
    .A3(_1156_),
    .B1(_1155_),
    .X(_1163_));
 sky130_fd_sc_hd__a21oi_1 _1723_ (.A1(_1118_),
    .A2(_1030_),
    .B1(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__and3_1 _1724_ (.A(_1118_),
    .B(_1030_),
    .C(_1163_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_1 _1725_ (.A(_1164_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__buf_2 _1726_ (.A(\m1.a[1] ),
    .X(_1167_));
 sky130_fd_sc_hd__nand2_1 _1727_ (.A(_1167_),
    .B(\m1.b[7] ),
    .Y(_1168_));
 sky130_fd_sc_hd__xor2_1 _1728_ (.A(_1166_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__nand2_1 _1729_ (.A(_1134_),
    .B(_1161_),
    .Y(_1170_));
 sky130_fd_sc_hd__xnor2_1 _1730_ (.A(_1160_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__and2b_1 _1731_ (.A_N(_1169_),
    .B(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__xor2_1 _1732_ (.A(_1123_),
    .B(_1137_),
    .X(_1173_));
 sky130_fd_sc_hd__o21ai_1 _1733_ (.A1(_1162_),
    .A2(_1172_),
    .B1(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__a31o_1 _1734_ (.A1(_1167_),
    .A2(_1029_),
    .A3(_1166_),
    .B1(_1165_),
    .X(_1175_));
 sky130_fd_sc_hd__or3_1 _1735_ (.A(_1162_),
    .B(_1172_),
    .C(_1173_),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _1736_ (.A(_1174_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__nand2_1 _1737_ (.A(_1175_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__xnor2_1 _1738_ (.A(_1121_),
    .B(_1142_),
    .Y(_1179_));
 sky130_fd_sc_hd__a21o_1 _1739_ (.A1(_1174_),
    .A2(_1178_),
    .B1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__xnor2_1 _1740_ (.A(_1175_),
    .B(_1177_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_1 _1741_ (.A(_1167_),
    .B(\m1.b[5] ),
    .Y(_1182_));
 sky130_fd_sc_hd__a22oi_1 _1742_ (.A1(\m1.a[2] ),
    .A2(_1038_),
    .B1(\m1.b[3] ),
    .B2(_1091_),
    .Y(_1183_));
 sky130_fd_sc_hd__and4_1 _1743_ (.A(\m1.a[3] ),
    .B(\m1.a[2] ),
    .C(\m1.b[4] ),
    .D(\m1.b[3] ),
    .X(_1184_));
 sky130_fd_sc_hd__nor2_1 _1744_ (.A(_1183_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__xnor2_1 _1745_ (.A(_1182_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__or3_1 _1746_ (.A(_1149_),
    .B(_1147_),
    .C(_1148_),
    .X(_1187_));
 sky130_fd_sc_hd__o21ai_1 _1747_ (.A1(_1149_),
    .A2(_1148_),
    .B1(_1147_),
    .Y(_1188_));
 sky130_fd_sc_hd__a22oi_2 _1748_ (.A1(\m1.a[4] ),
    .A2(\m1.b[1] ),
    .B1(\m1.b[0] ),
    .B2(\m1.a[5] ),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _1749_ (.A(\m1.a[3] ),
    .B(_1076_),
    .Y(_1190_));
 sky130_fd_sc_hd__and4_1 _1750_ (.A(\m1.a[5] ),
    .B(\m1.a[4] ),
    .C(\m1.b[1] ),
    .D(\m1.b[0] ),
    .X(_1191_));
 sky130_fd_sc_hd__o21bai_1 _1751_ (.A1(_1189_),
    .A2(_1190_),
    .B1_N(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__a21o_1 _1752_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__nand3_1 _1753_ (.A(_1187_),
    .B(_1192_),
    .C(_1188_),
    .Y(_1194_));
 sky130_fd_sc_hd__a21bo_1 _1754_ (.A1(_1186_),
    .A2(_1193_),
    .B1_N(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__a21o_1 _1755_ (.A1(_1152_),
    .A2(_1158_),
    .B1(_1157_),
    .X(_1196_));
 sky130_fd_sc_hd__nand3_1 _1756_ (.A(_1159_),
    .B(_1195_),
    .C(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__o21bai_1 _1757_ (.A1(_1182_),
    .A2(_1183_),
    .B1_N(_1184_),
    .Y(_1198_));
 sky130_fd_sc_hd__and2_1 _1758_ (.A(_1167_),
    .B(\m1.b[6] ),
    .X(_1199_));
 sky130_fd_sc_hd__nor2_1 _1759_ (.A(_1198_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__and2_1 _1760_ (.A(_1198_),
    .B(_1199_),
    .X(_1201_));
 sky130_fd_sc_hd__nor2_1 _1761_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__buf_2 _1762_ (.A(\m1.a[0] ),
    .X(_1203_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_1203_),
    .B(\m1.b[7] ),
    .Y(_1204_));
 sky130_fd_sc_hd__xnor2_1 _1764_ (.A(_1202_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__a21o_1 _1765_ (.A1(_1159_),
    .A2(_1196_),
    .B1(_1195_),
    .X(_1206_));
 sky130_fd_sc_hd__nand3_1 _1766_ (.A(_1197_),
    .B(_1205_),
    .C(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__and2_1 _1767_ (.A(_1197_),
    .B(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__xor2_1 _1768_ (.A(_1169_),
    .B(_1171_),
    .X(_1209_));
 sky130_fd_sc_hd__o21ba_1 _1769_ (.A1(_1200_),
    .A2(_1204_),
    .B1_N(_1201_),
    .X(_1210_));
 sky130_fd_sc_hd__xor2_1 _1770_ (.A(_1208_),
    .B(_1209_),
    .X(_1211_));
 sky130_fd_sc_hd__or2b_1 _1771_ (.A(_1210_),
    .B_N(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__o21ai_1 _1772_ (.A1(_1208_),
    .A2(_1209_),
    .B1(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__or2b_1 _1773_ (.A(_1181_),
    .B_N(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__nand3_1 _1774_ (.A(_1194_),
    .B(_1186_),
    .C(_1193_),
    .Y(_1215_));
 sky130_fd_sc_hd__a22o_1 _1775_ (.A1(\m1.a[1] ),
    .A2(\m1.b[4] ),
    .B1(\m1.b[3] ),
    .B2(\m1.a[2] ),
    .X(_1216_));
 sky130_fd_sc_hd__nand4_1 _1776_ (.A(_1118_),
    .B(\m1.a[1] ),
    .C(_1038_),
    .D(\m1.b[3] ),
    .Y(_1217_));
 sky130_fd_sc_hd__and2_1 _1777_ (.A(\m1.a[0] ),
    .B(\m1.b[5] ),
    .X(_1218_));
 sky130_fd_sc_hd__a21oi_1 _1778_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__and3_1 _1779_ (.A(_1218_),
    .B(_1216_),
    .C(_1217_),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_1 _1780_ (.A(_1219_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__or3_1 _1781_ (.A(_1191_),
    .B(_1189_),
    .C(_1190_),
    .X(_1222_));
 sky130_fd_sc_hd__o21ai_1 _1782_ (.A1(_1191_),
    .A2(_1189_),
    .B1(_1190_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(\m1.a[2] ),
    .B(_1076_),
    .Y(_1224_));
 sky130_fd_sc_hd__a22oi_2 _1784_ (.A1(\m1.a[3] ),
    .A2(_1077_),
    .B1(_1125_),
    .B2(\m1.a[4] ),
    .Y(_1225_));
 sky130_fd_sc_hd__and4_1 _1785_ (.A(\m1.a[4] ),
    .B(\m1.a[3] ),
    .C(\m1.b[1] ),
    .D(\m1.b[0] ),
    .X(_1226_));
 sky130_fd_sc_hd__o21bai_1 _1786_ (.A1(_1224_),
    .A2(_1225_),
    .B1_N(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__a21o_1 _1787_ (.A1(_1222_),
    .A2(_1223_),
    .B1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__nand3_1 _1788_ (.A(_1222_),
    .B(_1227_),
    .C(_1223_),
    .Y(_1229_));
 sky130_fd_sc_hd__a21bo_1 _1789_ (.A1(_1221_),
    .A2(_1228_),
    .B1_N(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__a21o_1 _1790_ (.A1(_1194_),
    .A2(_1193_),
    .B1(_1186_),
    .X(_1231_));
 sky130_fd_sc_hd__and3_1 _1791_ (.A(_1215_),
    .B(_1230_),
    .C(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__and4_1 _1792_ (.A(_1118_),
    .B(_1167_),
    .C(_1038_),
    .D(_1058_),
    .X(_1233_));
 sky130_fd_sc_hd__o211a_1 _1793_ (.A1(_1233_),
    .A2(_1220_),
    .B1(_1203_),
    .C1(\m1.b[6] ),
    .X(_1234_));
 sky130_fd_sc_hd__a211oi_1 _1794_ (.A1(_1203_),
    .A2(\m1.b[6] ),
    .B1(_1233_),
    .C1(_1220_),
    .Y(_1235_));
 sky130_fd_sc_hd__or2_1 _1795_ (.A(_1234_),
    .B(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__a21oi_1 _1796_ (.A1(_1215_),
    .A2(_1231_),
    .B1(_1230_),
    .Y(_1237_));
 sky130_fd_sc_hd__nor3_1 _1797_ (.A(_1232_),
    .B(_1236_),
    .C(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__a21o_1 _1798_ (.A1(_1197_),
    .A2(_1206_),
    .B1(_1205_),
    .X(_0260_));
 sky130_fd_sc_hd__o211a_1 _1799_ (.A1(_1232_),
    .A2(_1238_),
    .B1(_0260_),
    .C1(_1207_),
    .X(_0261_));
 sky130_fd_sc_hd__a211oi_1 _1800_ (.A1(_1207_),
    .A2(_0260_),
    .B1(_1238_),
    .C1(_1232_),
    .Y(_0262_));
 sky130_fd_sc_hd__or3b_1 _1801_ (.A(_0261_),
    .B(_0262_),
    .C_N(_1234_),
    .X(_0263_));
 sky130_fd_sc_hd__or2b_1 _1802_ (.A(_0261_),
    .B_N(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__xnor2_1 _1803_ (.A(_1210_),
    .B(_1211_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _1804_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3_1 _1805_ (.A(_1229_),
    .B(_1221_),
    .C(_1228_),
    .Y(_0267_));
 sky130_fd_sc_hd__a22o_1 _1806_ (.A1(\m1.a[0] ),
    .A2(_1038_),
    .B1(_1058_),
    .B2(_1167_),
    .X(_0268_));
 sky130_fd_sc_hd__and4_1 _1807_ (.A(\m1.a[1] ),
    .B(\m1.a[0] ),
    .C(\m1.b[4] ),
    .D(\m1.b[3] ),
    .X(_0269_));
 sky130_fd_sc_hd__inv_2 _1808_ (.A(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__and2_1 _1809_ (.A(_0268_),
    .B(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__or3_1 _1810_ (.A(_1226_),
    .B(_1224_),
    .C(_1225_),
    .X(_0272_));
 sky130_fd_sc_hd__o21ai_1 _1811_ (.A1(_1226_),
    .A2(_1225_),
    .B1(_1224_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _1812_ (.A(_1167_),
    .B(_1076_),
    .Y(_0274_));
 sky130_fd_sc_hd__a22oi_1 _1813_ (.A1(_1118_),
    .A2(_1077_),
    .B1(_1125_),
    .B2(_1091_),
    .Y(_0275_));
 sky130_fd_sc_hd__and4_1 _1814_ (.A(\m1.a[3] ),
    .B(\m1.a[2] ),
    .C(\m1.b[1] ),
    .D(\m1.b[0] ),
    .X(_0276_));
 sky130_fd_sc_hd__o21bai_1 _1815_ (.A1(_0274_),
    .A2(_0275_),
    .B1_N(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21o_1 _1816_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__and3_1 _1817_ (.A(_0272_),
    .B(_0277_),
    .C(_0273_),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _1818_ (.A1(_0271_),
    .A2(_0278_),
    .B1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _1819_ (.A1(_1229_),
    .A2(_1228_),
    .B1(_1221_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _1820_ (.A(_0267_),
    .B(_0280_),
    .C(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__a21oi_1 _1821_ (.A1(_0267_),
    .A2(_0281_),
    .B1(_0280_),
    .Y(_0283_));
 sky130_fd_sc_hd__nor3_1 _1822_ (.A(_0270_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _1823_ (.A1(_1232_),
    .A2(_1237_),
    .B1(_1236_),
    .Y(_0285_));
 sky130_fd_sc_hd__or3_1 _1824_ (.A(_1232_),
    .B(_1236_),
    .C(_1237_),
    .X(_0286_));
 sky130_fd_sc_hd__o211a_1 _1825_ (.A1(_0282_),
    .A2(_0284_),
    .B1(_0285_),
    .C1(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__o21bai_1 _1826_ (.A1(_0261_),
    .A2(_0262_),
    .B1_N(_1234_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand3_1 _1827_ (.A(_0263_),
    .B(_0287_),
    .C(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__and3_1 _1828_ (.A(_0263_),
    .B(_0287_),
    .C(_0288_),
    .X(_0290_));
 sky130_fd_sc_hd__a21oi_1 _1829_ (.A1(_0263_),
    .A2(_0288_),
    .B1(_0287_),
    .Y(_0291_));
 sky130_fd_sc_hd__a211oi_1 _1830_ (.A1(_0286_),
    .A2(_0285_),
    .B1(_0284_),
    .C1(_0282_),
    .Y(_0292_));
 sky130_fd_sc_hd__and4_1 _1831_ (.A(\m1.a[2] ),
    .B(\m1.a[1] ),
    .C(\m1.b[1] ),
    .D(_1125_),
    .X(_0293_));
 sky130_fd_sc_hd__a22oi_1 _1832_ (.A1(\m1.a[1] ),
    .A2(_1077_),
    .B1(_1125_),
    .B2(_1118_),
    .Y(_0294_));
 sky130_fd_sc_hd__and4bb_1 _1833_ (.A_N(_0293_),
    .B_N(_0294_),
    .C(\m1.a[0] ),
    .D(_1076_),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_1 _1834_ (.A(_0293_),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__nor2_1 _1835_ (.A(_0276_),
    .B(_0275_),
    .Y(_0297_));
 sky130_fd_sc_hd__xnor2_1 _1836_ (.A(_0274_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__and2b_1 _1837_ (.A_N(_0296_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__xnor2_1 _1838_ (.A(_0296_),
    .B(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__and3_1 _1839_ (.A(_1203_),
    .B(_1058_),
    .C(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__and2b_1 _1840_ (.A_N(_0279_),
    .B(_0278_),
    .X(_0302_));
 sky130_fd_sc_hd__xor2_1 _1841_ (.A(_0271_),
    .B(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__o21ai_2 _1842_ (.A1(_0299_),
    .A2(_0301_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__o21a_1 _1843_ (.A1(_0282_),
    .A2(_0283_),
    .B1(_0270_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _1844_ (.A(_0284_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__o22a_1 _1845_ (.A1(_0287_),
    .A2(_0292_),
    .B1(_0304_),
    .B2(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__and4_1 _1846_ (.A(_1167_),
    .B(_1203_),
    .C(_1077_),
    .D(_1125_),
    .X(_0308_));
 sky130_fd_sc_hd__o2bb2a_1 _1847_ (.A1_N(_1203_),
    .A2_N(_1076_),
    .B1(_0293_),
    .B2(_0294_),
    .X(_0309_));
 sky130_fd_sc_hd__nor2_1 _1848_ (.A(_0295_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__and2_1 _1849_ (.A(_0308_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_1 _1850_ (.A(_1203_),
    .B(_1058_),
    .Y(_0312_));
 sky130_fd_sc_hd__xnor2_1 _1851_ (.A(_0312_),
    .B(_0300_),
    .Y(_0313_));
 sky130_fd_sc_hd__and2_1 _1852_ (.A(_0311_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__or3_1 _1853_ (.A(_0303_),
    .B(_0299_),
    .C(_0301_),
    .X(_0315_));
 sky130_fd_sc_hd__nand3_1 _1854_ (.A(_0304_),
    .B(_0314_),
    .C(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2_1 _1855_ (.A(_0306_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__nor4_1 _1856_ (.A(_0287_),
    .B(_0292_),
    .C(_0304_),
    .D(_0306_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21ba_1 _1857_ (.A1(_0307_),
    .A2(_0317_),
    .B1_N(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _1858_ (.A(_0290_),
    .B(_0291_),
    .C(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__xnor2_1 _1859_ (.A(_0264_),
    .B(_0265_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_1 _1860_ (.A1(_0289_),
    .A2(_0320_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__xor2_1 _1861_ (.A(_1213_),
    .B(_1181_),
    .X(_0323_));
 sky130_fd_sc_hd__a21o_1 _1862_ (.A1(_0266_),
    .A2(_0322_),
    .B1(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__nand3_1 _1863_ (.A(_1174_),
    .B(_1178_),
    .C(_1179_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _1864_ (.A(_1180_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__a21o_1 _1865_ (.A1(_1214_),
    .A2(_0324_),
    .B1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__xor2_1 _1866_ (.A(_1144_),
    .B(_1111_),
    .X(_0328_));
 sky130_fd_sc_hd__a21o_1 _1867_ (.A1(_1180_),
    .A2(_0327_),
    .B1(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nand3_1 _1868_ (.A(_1103_),
    .B(_1107_),
    .C(_1109_),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _1869_ (.A(_1110_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__a21o_1 _1870_ (.A1(_1145_),
    .A2(_0329_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nand3_1 _1871_ (.A(_1069_),
    .B(_1072_),
    .C(_1074_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _1872_ (.A(_1075_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21o_1 _1873_ (.A1(_1110_),
    .A2(_0332_),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__xnor2_1 _1874_ (.A(_1051_),
    .B(_1052_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _1875_ (.A1(_1075_),
    .A2(_0335_),
    .B1(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__or2_1 _1876_ (.A(_0993_),
    .B(\m1.multa_reg[15] ),
    .X(_0338_));
 sky130_fd_sc_hd__o31a_1 _1877_ (.A1(_0988_),
    .A2(_1053_),
    .A3(_0337_),
    .B1(_0338_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _1878_ (.A(_0336_),
    .B(_1075_),
    .C(_0335_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _1879_ (.A(_0988_),
    .B(\m1.multa_reg[14] ),
    .Y(_0340_));
 sky130_fd_sc_hd__o31ai_1 _1880_ (.A1(_0988_),
    .A2(_0337_),
    .A3(_0339_),
    .B1(_0340_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand3_1 _1881_ (.A(_0334_),
    .B(_1110_),
    .C(_0332_),
    .Y(_0341_));
 sky130_fd_sc_hd__and3_1 _1882_ (.A(_0993_),
    .B(_0335_),
    .C(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a21o_1 _1883_ (.A1(_0992_),
    .A2(\m1.multa_reg[13] ),
    .B1(_0342_),
    .X(_0241_));
 sky130_fd_sc_hd__nand3_1 _1884_ (.A(_0331_),
    .B(_1145_),
    .C(_0329_),
    .Y(_0343_));
 sky130_fd_sc_hd__and2_1 _1885_ (.A(_0991_),
    .B(\m1.multa_reg[12] ),
    .X(_0344_));
 sky130_fd_sc_hd__a31o_1 _1886_ (.A1(_0985_),
    .A2(_0332_),
    .A3(_0343_),
    .B1(_0344_),
    .X(_0240_));
 sky130_fd_sc_hd__nand3_1 _1887_ (.A(_0328_),
    .B(_1180_),
    .C(_0327_),
    .Y(_0345_));
 sky130_fd_sc_hd__and2_1 _1888_ (.A(_0991_),
    .B(\m1.multa_reg[11] ),
    .X(_0346_));
 sky130_fd_sc_hd__a31o_1 _1889_ (.A1(_0985_),
    .A2(_0329_),
    .A3(_0345_),
    .B1(_0346_),
    .X(_0239_));
 sky130_fd_sc_hd__nand3_1 _1890_ (.A(_0326_),
    .B(_1214_),
    .C(_0324_),
    .Y(_0347_));
 sky130_fd_sc_hd__and2_1 _1891_ (.A(_0991_),
    .B(\m1.multa_reg[10] ),
    .X(_0348_));
 sky130_fd_sc_hd__a31o_1 _1892_ (.A1(_0985_),
    .A2(_0327_),
    .A3(_0347_),
    .B1(_0348_),
    .X(_0238_));
 sky130_fd_sc_hd__nand3_1 _1893_ (.A(_0323_),
    .B(_0266_),
    .C(_0322_),
    .Y(_0349_));
 sky130_fd_sc_hd__and2_1 _1894_ (.A(_0987_),
    .B(\m1.multa_reg[9] ),
    .X(_0350_));
 sky130_fd_sc_hd__a31o_1 _1895_ (.A1(_0985_),
    .A2(_0324_),
    .A3(_0349_),
    .B1(_0350_),
    .X(_0237_));
 sky130_fd_sc_hd__nand3_1 _1896_ (.A(_0321_),
    .B(_0289_),
    .C(_0320_),
    .Y(_0351_));
 sky130_fd_sc_hd__and2_1 _1897_ (.A(_0987_),
    .B(\m1.multa_reg[8] ),
    .X(_0352_));
 sky130_fd_sc_hd__a31o_1 _1898_ (.A1(_0985_),
    .A2(_0322_),
    .A3(_0351_),
    .B1(_0352_),
    .X(_0236_));
 sky130_fd_sc_hd__o21ai_1 _1899_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0319_),
    .Y(_0353_));
 sky130_fd_sc_hd__and2_1 _1900_ (.A(_0987_),
    .B(\m1.multa_reg[7] ),
    .X(_0354_));
 sky130_fd_sc_hd__a31o_1 _1901_ (.A1(_0985_),
    .A2(_0320_),
    .A3(_0353_),
    .B1(_0354_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _1902_ (.A(_0318_),
    .B(_0307_),
    .X(_0355_));
 sky130_fd_sc_hd__xor2_1 _1903_ (.A(_0355_),
    .B(_0317_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _1904_ (.A0(\m1.multa_reg[6] ),
    .A1(_0356_),
    .S(_1012_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _1905_ (.A(_0357_),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _1906_ (.A(_0304_),
    .B(_0316_),
    .Y(_0358_));
 sky130_fd_sc_hd__xnor2_1 _1907_ (.A(_0306_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(\m1.multa_reg[5] ),
    .A1(_0359_),
    .S(_1012_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _1909_ (.A(_0360_),
    .X(_0233_));
 sky130_fd_sc_hd__a21o_1 _1910_ (.A1(_0304_),
    .A2(_0315_),
    .B1(_0314_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _1911_ (.A(_0987_),
    .B(\m1.multa_reg[4] ),
    .X(_0362_));
 sky130_fd_sc_hd__a31o_1 _1912_ (.A1(_0985_),
    .A2(_0316_),
    .A3(_0361_),
    .B1(_0362_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _1913_ (.A(_0311_),
    .B(_0313_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_1 _1914_ (.A(_0314_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(\m1.multa_reg[3] ),
    .A1(_0364_),
    .S(_1012_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _1916_ (.A(_0365_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _1917_ (.A(_0308_),
    .B(_0310_),
    .X(_0366_));
 sky130_fd_sc_hd__nor2_1 _1918_ (.A(_0991_),
    .B(_0311_),
    .Y(_0367_));
 sky130_fd_sc_hd__a22o_1 _1919_ (.A1(_0988_),
    .A2(\m1.multa_reg[2] ),
    .B1(_0366_),
    .B2(_0367_),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _1920_ (.A1(_1203_),
    .A2(_1077_),
    .B1(_1125_),
    .B2(_1167_),
    .X(_0368_));
 sky130_fd_sc_hd__and3b_1 _1921_ (.A_N(_0308_),
    .B(_0368_),
    .C(_0993_),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _1922_ (.A1(_0992_),
    .A2(\m1.multa_reg[1] ),
    .B1(_0369_),
    .X(_0229_));
 sky130_fd_sc_hd__and3_1 _1923_ (.A(_0993_),
    .B(_1203_),
    .C(_1125_),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _1924_ (.A1(_0992_),
    .A2(\m1.multa_reg[0] ),
    .B1(_0370_),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _1925_ (.A(\m2.multa_reg[15] ),
    .B(\m2.out[15] ),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _1926_ (.A(\m2.multa_reg[14] ),
    .B(\m2.out[14] ),
    .Y(_0372_));
 sky130_fd_sc_hd__or2_1 _1927_ (.A(\m2.multa_reg[13] ),
    .B(\m2.out[13] ),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_1 _1928_ (.A(\m2.multa_reg[12] ),
    .B(\m2.out[12] ),
    .Y(_0374_));
 sky130_fd_sc_hd__or2_1 _1929_ (.A(\m2.multa_reg[11] ),
    .B(\m2.out[11] ),
    .X(_0375_));
 sky130_fd_sc_hd__nor2_1 _1930_ (.A(\m2.multa_reg[10] ),
    .B(\m2.out[10] ),
    .Y(_0376_));
 sky130_fd_sc_hd__or2_1 _1931_ (.A(\m2.multa_reg[9] ),
    .B(\m2.out[9] ),
    .X(_0377_));
 sky130_fd_sc_hd__nor2_1 _1932_ (.A(\m2.multa_reg[8] ),
    .B(\m2.out[8] ),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _1933_ (.A(\m2.multa_reg[7] ),
    .B(\m2.out[7] ),
    .Y(_0379_));
 sky130_fd_sc_hd__nor2_1 _1934_ (.A(\m2.multa_reg[6] ),
    .B(\m2.out[6] ),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _1935_ (.A(\m2.multa_reg[5] ),
    .B(\m2.out[5] ),
    .Y(_0381_));
 sky130_fd_sc_hd__and2_1 _1936_ (.A(\m2.multa_reg[4] ),
    .B(\m2.out[4] ),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _1937_ (.A(\m2.multa_reg[4] ),
    .B(\m2.out[4] ),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_1 _1938_ (.A(_0382_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__or2_1 _1939_ (.A(\m2.multa_reg[3] ),
    .B(\m2.out[3] ),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _1940_ (.A(\m2.multa_reg[2] ),
    .B(\m2.out[2] ),
    .Y(_0386_));
 sky130_fd_sc_hd__nand2_1 _1941_ (.A(\m2.multa_reg[1] ),
    .B(\m2.out[1] ),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_1 _1942_ (.A(\m2.multa_reg[1] ),
    .B(\m2.out[1] ),
    .X(_0388_));
 sky130_fd_sc_hd__and4_1 _1943_ (.A(\m2.multa_reg[0] ),
    .B(\m2.out[0] ),
    .C(_0387_),
    .D(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__a21oi_1 _1944_ (.A1(\m2.multa_reg[1] ),
    .A2(\m2.out[1] ),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_1 _1945_ (.A(\m2.multa_reg[2] ),
    .B(\m2.out[2] ),
    .Y(_0391_));
 sky130_fd_sc_hd__o21ai_1 _1946_ (.A1(_0386_),
    .A2(_0390_),
    .B1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21o_1 _1947_ (.A1(\m2.multa_reg[3] ),
    .A2(\m2.out[3] ),
    .B1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__a31oi_2 _1948_ (.A1(_0384_),
    .A2(_0385_),
    .A3(_0393_),
    .B1(_0382_),
    .Y(_0394_));
 sky130_fd_sc_hd__and2_1 _1949_ (.A(\m2.multa_reg[5] ),
    .B(\m2.out[5] ),
    .X(_0395_));
 sky130_fd_sc_hd__o21ba_1 _1950_ (.A1(_0381_),
    .A2(_0394_),
    .B1_N(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _1951_ (.A(\m2.multa_reg[6] ),
    .B(\m2.out[6] ),
    .Y(_0397_));
 sky130_fd_sc_hd__o21a_1 _1952_ (.A1(_0380_),
    .A2(_0396_),
    .B1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _1953_ (.A(\m2.multa_reg[7] ),
    .B(\m2.out[7] ),
    .Y(_0399_));
 sky130_fd_sc_hd__o21a_1 _1954_ (.A1(_0379_),
    .A2(_0398_),
    .B1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(\m2.multa_reg[8] ),
    .B(\m2.out[8] ),
    .Y(_0401_));
 sky130_fd_sc_hd__o21ai_1 _1956_ (.A1(_0378_),
    .A2(_0400_),
    .B1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _1957_ (.A(\m2.multa_reg[9] ),
    .B(\m2.out[9] ),
    .Y(_0403_));
 sky130_fd_sc_hd__a21boi_1 _1958_ (.A1(_0377_),
    .A2(_0402_),
    .B1_N(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _1959_ (.A(\m2.multa_reg[10] ),
    .B(\m2.out[10] ),
    .Y(_0405_));
 sky130_fd_sc_hd__o21ai_1 _1960_ (.A1(_0376_),
    .A2(_0404_),
    .B1(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(\m2.multa_reg[11] ),
    .B(\m2.out[11] ),
    .Y(_0407_));
 sky130_fd_sc_hd__a21boi_1 _1962_ (.A1(_0375_),
    .A2(_0406_),
    .B1_N(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _1963_ (.A(\m2.multa_reg[12] ),
    .B(\m2.out[12] ),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ai_1 _1964_ (.A1(_0374_),
    .A2(_0408_),
    .B1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(\m2.multa_reg[13] ),
    .B(\m2.out[13] ),
    .Y(_0411_));
 sky130_fd_sc_hd__a21boi_1 _1966_ (.A1(_0373_),
    .A2(_0410_),
    .B1_N(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _1967_ (.A(\m2.multa_reg[14] ),
    .B(\m2.out[14] ),
    .Y(_0413_));
 sky130_fd_sc_hd__o21ai_1 _1968_ (.A1(_0372_),
    .A2(_0412_),
    .B1(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__or2_1 _1969_ (.A(\m2.multa_reg[15] ),
    .B(\m2.out[15] ),
    .X(_0415_));
 sky130_fd_sc_hd__o211a_1 _1970_ (.A1(_0371_),
    .A2(_0414_),
    .B1(_0415_),
    .C1(_0984_),
    .X(_0416_));
 sky130_fd_sc_hd__xor2_1 _1971_ (.A(\m2.out[16] ),
    .B(_0416_),
    .X(_0227_));
 sky130_fd_sc_hd__or2b_1 _1972_ (.A(_0371_),
    .B_N(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1973_ (.A0(\m2.multa_reg[15] ),
    .A1(_0414_),
    .S(_0984_),
    .X(_0418_));
 sky130_fd_sc_hd__xnor2_1 _1974_ (.A(_0417_),
    .B(_0418_),
    .Y(_0226_));
 sky130_fd_sc_hd__and2b_1 _1975_ (.A_N(_0372_),
    .B(_0413_),
    .X(_0419_));
 sky130_fd_sc_hd__xnor2_1 _1976_ (.A(_0412_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(\m2.out[14] ),
    .A1(_0420_),
    .S(_1012_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1978_ (.A(_0421_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _1979_ (.A(_0373_),
    .B(_0411_),
    .Y(_0422_));
 sky130_fd_sc_hd__xnor2_1 _1980_ (.A(_0410_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__mux2_1 _1981_ (.A0(\m2.out[13] ),
    .A1(_0423_),
    .S(_1012_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1982_ (.A(_0424_),
    .X(_0224_));
 sky130_fd_sc_hd__and2b_1 _1983_ (.A_N(_0374_),
    .B(_0409_),
    .X(_0425_));
 sky130_fd_sc_hd__xnor2_1 _1984_ (.A(_0408_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__mux2_1 _1985_ (.A0(\m2.out[12] ),
    .A1(_0426_),
    .S(_1012_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _1986_ (.A(_0427_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(_0375_),
    .B(_0407_),
    .Y(_0428_));
 sky130_fd_sc_hd__xnor2_1 _1988_ (.A(_0406_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__mux2_1 _1989_ (.A0(\m2.out[11] ),
    .A1(_0429_),
    .S(_1012_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1990_ (.A(_0430_),
    .X(_0222_));
 sky130_fd_sc_hd__and2b_1 _1991_ (.A_N(_0376_),
    .B(_0405_),
    .X(_0431_));
 sky130_fd_sc_hd__xnor2_1 _1992_ (.A(_0404_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__buf_4 _1993_ (.A(net1),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(\m2.out[10] ),
    .A1(_0432_),
    .S(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1995_ (.A(_0434_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _1996_ (.A(_0377_),
    .B(_0403_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _1997_ (.A(_0402_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_1 _1998_ (.A0(\m2.out[9] ),
    .A1(_0436_),
    .S(_0433_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1999_ (.A(_0437_),
    .X(_0220_));
 sky130_fd_sc_hd__and2b_1 _2000_ (.A_N(_0378_),
    .B(_0401_),
    .X(_0438_));
 sky130_fd_sc_hd__xnor2_1 _2001_ (.A(_0400_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(\m2.out[8] ),
    .A1(_0439_),
    .S(_0433_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _2003_ (.A(_0440_),
    .X(_0219_));
 sky130_fd_sc_hd__and2b_1 _2004_ (.A_N(_0379_),
    .B(_0399_),
    .X(_0441_));
 sky130_fd_sc_hd__xnor2_1 _2005_ (.A(_0398_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__mux2_1 _2006_ (.A0(\m2.out[7] ),
    .A1(_0442_),
    .S(_0433_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _2007_ (.A(_0443_),
    .X(_0218_));
 sky130_fd_sc_hd__and2b_1 _2008_ (.A_N(_0380_),
    .B(_0397_),
    .X(_0444_));
 sky130_fd_sc_hd__xnor2_1 _2009_ (.A(_0396_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__mux2_1 _2010_ (.A0(\m2.out[6] ),
    .A1(_0445_),
    .S(_0433_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _2011_ (.A(_0446_),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _2012_ (.A(_0395_),
    .B(_0381_),
    .Y(_0447_));
 sky130_fd_sc_hd__xnor2_1 _2013_ (.A(_0447_),
    .B(_0394_),
    .Y(_0448_));
 sky130_fd_sc_hd__mux2_1 _2014_ (.A0(\m2.out[5] ),
    .A1(_0448_),
    .S(_0433_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _2015_ (.A(_0449_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_1 _2016_ (.A(_0385_),
    .B(_0393_),
    .Y(_0450_));
 sky130_fd_sc_hd__xnor2_1 _2017_ (.A(_0384_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__mux2_1 _2018_ (.A0(\m2.out[4] ),
    .A1(_0451_),
    .S(_0433_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _2019_ (.A(_0452_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _2020_ (.A(\m2.multa_reg[3] ),
    .B(\m2.out[3] ),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(_0385_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__xnor2_1 _2022_ (.A(_0392_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(\m2.out[3] ),
    .A1(_0455_),
    .S(_0433_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _2024_ (.A(_0456_),
    .X(_0214_));
 sky130_fd_sc_hd__and2b_1 _2025_ (.A_N(_0386_),
    .B(_0391_),
    .X(_0457_));
 sky130_fd_sc_hd__xnor2_1 _2026_ (.A(_0390_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(\m2.out[2] ),
    .A1(_0458_),
    .S(_0433_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _2028_ (.A(_0459_),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _2029_ (.A1(\m2.multa_reg[0] ),
    .A2(\m2.out[0] ),
    .B1(_0387_),
    .B2(_0388_),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _2030_ (.A(_0991_),
    .B(_0389_),
    .Y(_0461_));
 sky130_fd_sc_hd__a22o_1 _2031_ (.A1(_0988_),
    .A2(\m2.out[1] ),
    .B1(_0460_),
    .B2(_0461_),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(_0993_),
    .B(\m2.multa_reg[0] ),
    .Y(_0462_));
 sky130_fd_sc_hd__xnor2_1 _2033_ (.A(\m2.out[0] ),
    .B(_0462_),
    .Y(_0211_));
 sky130_fd_sc_hd__mux2_1 _2034_ (.A0(_0696_),
    .A1(\I3.out[7] ),
    .S(_0433_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _2035_ (.A(_0463_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_4 _2036_ (.A(net1),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2037_ (.A0(_0697_),
    .A1(\I3.out[6] ),
    .S(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _2038_ (.A(_0465_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(_0703_),
    .A1(\I3.out[5] ),
    .S(_0464_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _2040_ (.A(_0466_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2041_ (.A0(_0730_),
    .A1(\I3.out[4] ),
    .S(_0464_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _2042_ (.A(_0467_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _2043_ (.A0(_0747_),
    .A1(\I3.out[3] ),
    .S(_0464_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _2044_ (.A(_0468_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2045_ (.A0(_0783_),
    .A1(\I3.out[2] ),
    .S(_0464_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _2046_ (.A(_0469_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2047_ (.A0(_0813_),
    .A1(\I3.out[1] ),
    .S(_0464_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _2048_ (.A(_0470_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2049_ (.A0(_0869_),
    .A1(\I3.out[0] ),
    .S(_0464_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _2050_ (.A(_0471_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(_0698_),
    .A1(\I4.out[7] ),
    .S(_0464_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(_0472_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(_0699_),
    .A1(\I4.out[6] ),
    .S(_0464_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _2054_ (.A(_0473_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2055_ (.A0(_0702_),
    .A1(\I4.out[5] ),
    .S(_0464_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _2056_ (.A(_0474_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_4 _2057_ (.A(net1),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _2058_ (.A0(_0706_),
    .A1(\I4.out[4] ),
    .S(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _2059_ (.A(_0476_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(_0723_),
    .A1(\I4.out[3] ),
    .S(_0475_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _2061_ (.A(_0477_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(_0752_),
    .A1(\I4.out[2] ),
    .S(_0475_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _2063_ (.A(_0478_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2064_ (.A0(_0753_),
    .A1(\I4.out[1] ),
    .S(_0475_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _2065_ (.A(_0479_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(_0790_),
    .A1(\I4.out[0] ),
    .S(_0475_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _2067_ (.A(_0480_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_1 _2068_ (.A(\m1.multa_reg[15] ),
    .B(\m1.out[15] ),
    .X(_0481_));
 sky130_fd_sc_hd__nor2_1 _2069_ (.A(\m1.multa_reg[14] ),
    .B(\m1.out[14] ),
    .Y(_0482_));
 sky130_fd_sc_hd__or2_1 _2070_ (.A(\m1.multa_reg[13] ),
    .B(\m1.out[13] ),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_1 _2071_ (.A(\m1.multa_reg[12] ),
    .B(\m1.out[12] ),
    .Y(_0484_));
 sky130_fd_sc_hd__or2_1 _2072_ (.A(\m1.multa_reg[11] ),
    .B(\m1.out[11] ),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(\m1.multa_reg[10] ),
    .B(\m1.out[10] ),
    .Y(_0486_));
 sky130_fd_sc_hd__or2_1 _2074_ (.A(\m1.multa_reg[9] ),
    .B(\m1.out[9] ),
    .X(_0487_));
 sky130_fd_sc_hd__nor2_1 _2075_ (.A(\m1.multa_reg[8] ),
    .B(\m1.out[8] ),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _2076_ (.A(\m1.multa_reg[7] ),
    .B(\m1.out[7] ),
    .Y(_0489_));
 sky130_fd_sc_hd__nor2_1 _2077_ (.A(\m1.multa_reg[6] ),
    .B(\m1.out[6] ),
    .Y(_0490_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(\m1.multa_reg[5] ),
    .B(\m1.out[5] ),
    .Y(_0491_));
 sky130_fd_sc_hd__and2_1 _2079_ (.A(\m1.multa_reg[4] ),
    .B(\m1.out[4] ),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _2080_ (.A(\m1.multa_reg[4] ),
    .B(\m1.out[4] ),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(_0492_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_1 _2082_ (.A(\m1.multa_reg[3] ),
    .B(\m1.out[3] ),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_1 _2083_ (.A(\m1.multa_reg[2] ),
    .B(\m1.out[2] ),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _2084_ (.A(\m1.multa_reg[1] ),
    .B(\m1.out[1] ),
    .Y(_0497_));
 sky130_fd_sc_hd__or2_1 _2085_ (.A(\m1.multa_reg[1] ),
    .B(\m1.out[1] ),
    .X(_0498_));
 sky130_fd_sc_hd__and4_1 _2086_ (.A(\m1.multa_reg[0] ),
    .B(\m1.out[0] ),
    .C(_0497_),
    .D(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a21oi_1 _2087_ (.A1(\m1.multa_reg[1] ),
    .A2(\m1.out[1] ),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _2088_ (.A(\m1.multa_reg[2] ),
    .B(\m1.out[2] ),
    .Y(_0501_));
 sky130_fd_sc_hd__o21ai_1 _2089_ (.A1(_0496_),
    .A2(_0500_),
    .B1(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21o_1 _2090_ (.A1(\m1.multa_reg[3] ),
    .A2(\m1.out[3] ),
    .B1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a31oi_2 _2091_ (.A1(_0494_),
    .A2(_0495_),
    .A3(_0503_),
    .B1(_0492_),
    .Y(_0504_));
 sky130_fd_sc_hd__and2_1 _2092_ (.A(\m1.multa_reg[5] ),
    .B(\m1.out[5] ),
    .X(_0505_));
 sky130_fd_sc_hd__o21ba_1 _2093_ (.A1(_0491_),
    .A2(_0504_),
    .B1_N(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _2094_ (.A(\m1.multa_reg[6] ),
    .B(\m1.out[6] ),
    .Y(_0507_));
 sky130_fd_sc_hd__o21a_1 _2095_ (.A1(_0490_),
    .A2(_0506_),
    .B1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nand2_1 _2096_ (.A(\m1.multa_reg[7] ),
    .B(\m1.out[7] ),
    .Y(_0509_));
 sky130_fd_sc_hd__o21a_1 _2097_ (.A1(_0489_),
    .A2(_0508_),
    .B1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _2098_ (.A(\m1.multa_reg[8] ),
    .B(\m1.out[8] ),
    .Y(_0511_));
 sky130_fd_sc_hd__o21ai_1 _2099_ (.A1(_0488_),
    .A2(_0510_),
    .B1(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand2_1 _2100_ (.A(\m1.multa_reg[9] ),
    .B(\m1.out[9] ),
    .Y(_0513_));
 sky130_fd_sc_hd__a21boi_1 _2101_ (.A1(_0487_),
    .A2(_0512_),
    .B1_N(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _2102_ (.A(\m1.multa_reg[10] ),
    .B(\m1.out[10] ),
    .Y(_0515_));
 sky130_fd_sc_hd__o21ai_1 _2103_ (.A1(_0486_),
    .A2(_0514_),
    .B1(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _2104_ (.A(\m1.multa_reg[11] ),
    .B(\m1.out[11] ),
    .Y(_0517_));
 sky130_fd_sc_hd__a21boi_1 _2105_ (.A1(_0485_),
    .A2(_0516_),
    .B1_N(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(\m1.multa_reg[12] ),
    .B(\m1.out[12] ),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_1 _2107_ (.A1(_0484_),
    .A2(_0518_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _2108_ (.A(\m1.multa_reg[13] ),
    .B(\m1.out[13] ),
    .Y(_0521_));
 sky130_fd_sc_hd__a21boi_1 _2109_ (.A1(_0483_),
    .A2(_0520_),
    .B1_N(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _2110_ (.A(\m1.multa_reg[14] ),
    .B(\m1.out[14] ),
    .Y(_0523_));
 sky130_fd_sc_hd__o21ai_1 _2111_ (.A1(_0482_),
    .A2(_0522_),
    .B1(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _2112_ (.A(\m1.multa_reg[15] ),
    .B(\m1.out[15] ),
    .X(_0525_));
 sky130_fd_sc_hd__o211a_1 _2113_ (.A1(_0481_),
    .A2(_0524_),
    .B1(_0525_),
    .C1(_0984_),
    .X(_0526_));
 sky130_fd_sc_hd__xor2_1 _2114_ (.A(\m1.out[16] ),
    .B(_0526_),
    .X(_0194_));
 sky130_fd_sc_hd__or2b_1 _2115_ (.A(_0481_),
    .B_N(_0525_),
    .X(_0527_));
 sky130_fd_sc_hd__xnor2_1 _2116_ (.A(_0524_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(\m1.out[15] ),
    .A1(_0528_),
    .S(_0475_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _2118_ (.A(_0529_),
    .X(_0193_));
 sky130_fd_sc_hd__and2b_1 _2119_ (.A_N(_0482_),
    .B(_0523_),
    .X(_0530_));
 sky130_fd_sc_hd__xnor2_1 _2120_ (.A(_0522_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(\m1.out[14] ),
    .A1(_0531_),
    .S(_0475_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _2122_ (.A(_0532_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _2123_ (.A(_0483_),
    .B(_0521_),
    .Y(_0533_));
 sky130_fd_sc_hd__xnor2_1 _2124_ (.A(_0520_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__mux2_1 _2125_ (.A0(\m1.out[13] ),
    .A1(_0534_),
    .S(_0475_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _2126_ (.A(_0535_),
    .X(_0191_));
 sky130_fd_sc_hd__and2b_1 _2127_ (.A_N(_0484_),
    .B(_0519_),
    .X(_0536_));
 sky130_fd_sc_hd__xnor2_1 _2128_ (.A(_0518_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__mux2_1 _2129_ (.A0(\m1.out[12] ),
    .A1(_0537_),
    .S(_0475_),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _2130_ (.A(_0538_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_1 _2131_ (.A(_0485_),
    .B(_0517_),
    .Y(_0539_));
 sky130_fd_sc_hd__xnor2_1 _2132_ (.A(_0516_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(\m1.out[11] ),
    .A1(_0540_),
    .S(_0475_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _2134_ (.A(_0541_),
    .X(_0189_));
 sky130_fd_sc_hd__and2b_1 _2135_ (.A_N(_0486_),
    .B(_0515_),
    .X(_0542_));
 sky130_fd_sc_hd__xnor2_1 _2136_ (.A(_0514_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__buf_4 _2137_ (.A(net1),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(\m1.out[10] ),
    .A1(_0543_),
    .S(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__clkbuf_1 _2139_ (.A(_0545_),
    .X(_0188_));
 sky130_fd_sc_hd__nand2_1 _2140_ (.A(_0487_),
    .B(_0513_),
    .Y(_0546_));
 sky130_fd_sc_hd__xnor2_1 _2141_ (.A(_0512_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(\m1.out[9] ),
    .A1(_0547_),
    .S(_0544_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _2143_ (.A(_0548_),
    .X(_0187_));
 sky130_fd_sc_hd__and2b_1 _2144_ (.A_N(_0488_),
    .B(_0511_),
    .X(_0549_));
 sky130_fd_sc_hd__xnor2_1 _2145_ (.A(_0510_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__mux2_1 _2146_ (.A0(\m1.out[8] ),
    .A1(_0550_),
    .S(_0544_),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(_0551_),
    .X(_0186_));
 sky130_fd_sc_hd__and2b_1 _2148_ (.A_N(_0489_),
    .B(_0509_),
    .X(_0552_));
 sky130_fd_sc_hd__xnor2_1 _2149_ (.A(_0508_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\m1.out[7] ),
    .A1(_0553_),
    .S(_0544_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _2151_ (.A(_0554_),
    .X(_0185_));
 sky130_fd_sc_hd__and2b_1 _2152_ (.A_N(_0490_),
    .B(_0507_),
    .X(_0555_));
 sky130_fd_sc_hd__xnor2_1 _2153_ (.A(_0506_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__mux2_1 _2154_ (.A0(\m1.out[6] ),
    .A1(_0556_),
    .S(_0544_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _2155_ (.A(_0557_),
    .X(_0184_));
 sky130_fd_sc_hd__nor2_1 _2156_ (.A(_0505_),
    .B(_0491_),
    .Y(_0558_));
 sky130_fd_sc_hd__xnor2_1 _2157_ (.A(_0558_),
    .B(_0504_),
    .Y(_0559_));
 sky130_fd_sc_hd__mux2_1 _2158_ (.A0(\m1.out[5] ),
    .A1(_0559_),
    .S(_0544_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _2159_ (.A(_0560_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _2160_ (.A(_0495_),
    .B(_0503_),
    .Y(_0561_));
 sky130_fd_sc_hd__xnor2_1 _2161_ (.A(_0494_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2_1 _2162_ (.A0(\m1.out[4] ),
    .A1(_0562_),
    .S(_0544_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _2163_ (.A(_0563_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _2164_ (.A(\m1.multa_reg[3] ),
    .B(\m1.out[3] ),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _2165_ (.A(_0495_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__xnor2_1 _2166_ (.A(_0502_),
    .B(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(\m1.out[3] ),
    .A1(_0566_),
    .S(_0544_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _2168_ (.A(_0567_),
    .X(_0181_));
 sky130_fd_sc_hd__and2b_1 _2169_ (.A_N(_0496_),
    .B(_0501_),
    .X(_0568_));
 sky130_fd_sc_hd__xnor2_1 _2170_ (.A(_0500_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__mux2_1 _2171_ (.A0(\m1.out[2] ),
    .A1(_0569_),
    .S(_0544_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _2172_ (.A(_0570_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _2173_ (.A1(\m1.multa_reg[0] ),
    .A2(\m1.out[0] ),
    .B1(_0497_),
    .B2(_0498_),
    .X(_0571_));
 sky130_fd_sc_hd__nor2_1 _2174_ (.A(_0991_),
    .B(_0499_),
    .Y(_0572_));
 sky130_fd_sc_hd__a22o_1 _2175_ (.A1(_0988_),
    .A2(\m1.out[1] ),
    .B1(_0571_),
    .B2(_0572_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _2176_ (.A(_0993_),
    .B(\m1.multa_reg[0] ),
    .Y(_0573_));
 sky130_fd_sc_hd__xnor2_1 _2177_ (.A(\m1.out[0] ),
    .B(_0573_),
    .Y(_0178_));
 sky130_fd_sc_hd__mux2_1 _2178_ (.A0(_1027_),
    .A1(\I1.out[7] ),
    .S(_0544_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _2179_ (.A(_0574_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_4 _2180_ (.A(net1),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _2181_ (.A0(_1028_),
    .A1(\I1.out[6] ),
    .S(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _2182_ (.A(_0576_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2183_ (.A0(_1035_),
    .A1(\I1.out[5] ),
    .S(_0575_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _2184_ (.A(_0577_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2185_ (.A0(_1057_),
    .A1(\I1.out[4] ),
    .S(_0575_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _2186_ (.A(_0578_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2187_ (.A0(_1091_),
    .A1(\I1.out[3] ),
    .S(_0575_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _2188_ (.A(_0579_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2189_ (.A0(_1118_),
    .A1(\I1.out[2] ),
    .S(_0575_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _2190_ (.A(_0580_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2191_ (.A0(_1167_),
    .A1(\I1.out[1] ),
    .S(_0575_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _2192_ (.A(_0581_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(_1203_),
    .A1(\I1.out[0] ),
    .S(_0575_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_1 _2194_ (.A(_0582_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2195_ (.A0(_1029_),
    .A1(\I2.out[7] ),
    .S(_0575_),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _2196_ (.A(_0583_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(_1030_),
    .A1(\I2.out[6] ),
    .S(_0575_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _2198_ (.A(_0584_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(_1034_),
    .A1(\I2.out[5] ),
    .S(_0575_),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _2200_ (.A(_0585_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(_1038_),
    .A1(\I2.out[4] ),
    .S(_0984_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_1 _2202_ (.A(_0586_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(_1058_),
    .A1(\I2.out[3] ),
    .S(_0984_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _2204_ (.A(_0587_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2205_ (.A0(_1076_),
    .A1(\I2.out[2] ),
    .S(_0984_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_1 _2206_ (.A(_0588_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(_1077_),
    .A1(\I2.out[1] ),
    .S(_0984_),
    .X(_0589_));
 sky130_fd_sc_hd__clkbuf_1 _2208_ (.A(_0589_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(_1125_),
    .A1(\I2.out[0] ),
    .S(_0984_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_1 _2210_ (.A(_0590_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_2 _2211_ (.A(net10),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _2212_ (.A0(\P1.qq[9] ),
    .A1(\P1.in[1] ),
    .S(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_1 _2213_ (.A(_0592_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(\P1.qq[10] ),
    .A1(\P1.in[2] ),
    .S(_0591_),
    .X(_0593_));
 sky130_fd_sc_hd__clkbuf_1 _2215_ (.A(_0593_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(\P1.qq[11] ),
    .A1(\P1.in[3] ),
    .S(net10),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_1 _2217_ (.A(_0594_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2218_ (.A0(\P1.qq[12] ),
    .A1(\P1.in[4] ),
    .S(net10),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_1 _2219_ (.A(_0595_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(\P1.qq[13] ),
    .A1(\P1.in[5] ),
    .S(net10),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_1 _2221_ (.A(_0596_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(\P1.qq[14] ),
    .A1(\P1.in[6] ),
    .S(net10),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_1 _2223_ (.A(_0597_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(\P1.qq[15] ),
    .A1(\P1.in[7] ),
    .S(net10),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_1 _2225_ (.A(_0598_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _2226_ (.A(_0591_),
    .B(\P1.in[8] ),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(_0599_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _2228_ (.A(_0591_),
    .B(\P1.in[9] ),
    .X(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(_0600_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _2230_ (.A(_0591_),
    .B(\P1.in[10] ),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_0601_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _2232_ (.A(_0591_),
    .B(\P1.in[11] ),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_0602_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _2234_ (.A(_0591_),
    .B(\P1.in[12] ),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_0603_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _2236_ (.A(_0591_),
    .B(\P1.in[13] ),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(_0604_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _2238_ (.A(_0591_),
    .B(\P1.in[14] ),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_1 _2239_ (.A(_0605_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _2240_ (.A(_0591_),
    .B(\P1.in[15] ),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _2241_ (.A(_0606_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_2 _2242_ (.A(\A1.x[7] ),
    .X(_0607_));
 sky130_fd_sc_hd__inv_2 _2243_ (.A(net15),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_1 _2244_ (.A(_0607_),
    .B(_0016_),
    .Y(_0608_));
 sky130_fd_sc_hd__o21a_1 _2245_ (.A1(\A1.x[1] ),
    .A2(\A1.x[0] ),
    .B1(\A1.x[7] ),
    .X(_0609_));
 sky130_fd_sc_hd__a21o_1 _2246_ (.A1(\A1.x[2] ),
    .A2(\A1.x[7] ),
    .B1(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__xnor2_4 _2247_ (.A(\A1.x[3] ),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__xnor2_4 _2248_ (.A(\A1.x[2] ),
    .B(_0609_),
    .Y(_0612_));
 sky130_fd_sc_hd__or2b_1 _2249_ (.A(_0611_),
    .B_N(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_1 _2250_ (.A(_0608_),
    .B(_0613_),
    .Y(net17));
 sky130_fd_sc_hd__or4_1 _2251_ (.A(\A1.x[2] ),
    .B(\A1.x[1] ),
    .C(\A1.x[0] ),
    .D(\A1.x[3] ),
    .X(_0614_));
 sky130_fd_sc_hd__nand2_1 _2252_ (.A(\A1.x[7] ),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__xnor2_2 _2253_ (.A(\A1.x[4] ),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _2254_ (.A(_0611_),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__or2_1 _2255_ (.A(_0611_),
    .B(_0616_),
    .X(_0618_));
 sky130_fd_sc_hd__and2_1 _2256_ (.A(_0617_),
    .B(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _2257_ (.A(_0612_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__or2_1 _2258_ (.A(_0607_),
    .B(_0613_),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_0620_),
    .A2(_0621_),
    .B1(_0608_),
    .Y(net18));
 sky130_fd_sc_hd__inv_2 _2260_ (.A(_0607_),
    .Y(_0622_));
 sky130_fd_sc_hd__o21ai_2 _2261_ (.A1(\A1.x[4] ),
    .A2(_0614_),
    .B1(_0607_),
    .Y(_0623_));
 sky130_fd_sc_hd__xnor2_4 _2262_ (.A(\A1.x[5] ),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__or2_1 _2263_ (.A(_0616_),
    .B(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_1 _2264_ (.A(_0616_),
    .B(_0624_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _2265_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__mux2_1 _2266_ (.A0(_0627_),
    .A1(_0617_),
    .S(_0612_),
    .X(_0628_));
 sky130_fd_sc_hd__buf_4 _2267_ (.A(net15),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _2268_ (.A(_0620_),
    .B(_0627_),
    .Y(_0630_));
 sky130_fd_sc_hd__and3_1 _2269_ (.A(_0613_),
    .B(_0620_),
    .C(_0628_),
    .X(_0631_));
 sky130_fd_sc_hd__or4_1 _2270_ (.A(_0607_),
    .B(_0629_),
    .C(_0630_),
    .D(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__o21ai_1 _2271_ (.A1(_0622_),
    .A2(_0628_),
    .B1(_0632_),
    .Y(net19));
 sky130_fd_sc_hd__or2_1 _2272_ (.A(_0611_),
    .B(_0627_),
    .X(_0633_));
 sky130_fd_sc_hd__o31a_2 _2273_ (.A1(\A1.x[4] ),
    .A2(\A1.x[5] ),
    .A3(_0614_),
    .B1(\A1.x[7] ),
    .X(_0634_));
 sky130_fd_sc_hd__xor2_2 _2274_ (.A(\A1.x[6] ),
    .B(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or2_1 _2275_ (.A(_0612_),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_2 _2276_ (.A(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0626_),
    .A2(_0635_),
    .B1(_0612_),
    .Y(_0638_));
 sky130_fd_sc_hd__o21ai_1 _2278_ (.A1(_0626_),
    .A2(_0637_),
    .B1(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__xnor2_1 _2279_ (.A(_0633_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__and2_1 _2280_ (.A(_0631_),
    .B(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__nor2_1 _2281_ (.A(_0631_),
    .B(_0640_),
    .Y(_0642_));
 sky130_fd_sc_hd__or4_1 _2282_ (.A(_0607_),
    .B(net15),
    .C(_0641_),
    .D(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__o21ai_1 _2283_ (.A1(_0622_),
    .A2(_0640_),
    .B1(_0643_),
    .Y(net20));
 sky130_fd_sc_hd__or2_1 _2284_ (.A(_0611_),
    .B(_0635_),
    .X(_0644_));
 sky130_fd_sc_hd__or2_1 _2285_ (.A(_0619_),
    .B(_0635_),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_1 _2286_ (.A(_0637_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _2287_ (.A(_0620_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__and2b_1 _2288_ (.A_N(_0616_),
    .B(_0624_),
    .X(_0648_));
 sky130_fd_sc_hd__xnor2_1 _2289_ (.A(_0645_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__xor2_1 _2290_ (.A(_0647_),
    .B(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__xor2_1 _2291_ (.A(_0644_),
    .B(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _2292_ (.A(_0616_),
    .B(_0624_),
    .Y(_0652_));
 sky130_fd_sc_hd__a211o_1 _2293_ (.A1(_0626_),
    .A2(_0637_),
    .B1(_0611_),
    .C1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__xnor2_1 _2294_ (.A(_0651_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__o21ai_1 _2295_ (.A1(_0626_),
    .A2(_0637_),
    .B1(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and2_1 _2296_ (.A(_0641_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _2297_ (.A(_0607_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__o21a_1 _2298_ (.A1(_0641_),
    .A2(_0655_),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a2bb2o_1 _2299_ (.A1_N(_0622_),
    .A2_N(_0655_),
    .B1(_0658_),
    .B2(_0016_),
    .X(net21));
 sky130_fd_sc_hd__and3_1 _2300_ (.A(_0616_),
    .B(_0624_),
    .C(_0645_),
    .X(_0659_));
 sky130_fd_sc_hd__xnor2_2 _2301_ (.A(\A1.x[6] ),
    .B(_0634_),
    .Y(_0660_));
 sky130_fd_sc_hd__o2111a_1 _2302_ (.A1(_0612_),
    .A2(_0616_),
    .B1(_0617_),
    .C1(_0660_),
    .D1(_0613_),
    .X(_0661_));
 sky130_fd_sc_hd__a31oi_1 _2303_ (.A1(_0620_),
    .A2(_0646_),
    .A3(_0649_),
    .B1(_0659_),
    .Y(_0662_));
 sky130_fd_sc_hd__o32a_1 _2304_ (.A1(_0644_),
    .A2(_0659_),
    .A3(_0650_),
    .B1(_0661_),
    .B2(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__xnor2_1 _2305_ (.A(_0611_),
    .B(_0612_),
    .Y(_0664_));
 sky130_fd_sc_hd__xnor2_1 _2306_ (.A(_0624_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__a21oi_1 _2307_ (.A1(_0625_),
    .A2(_0633_),
    .B1(_0635_),
    .Y(_0666_));
 sky130_fd_sc_hd__a21oi_1 _2308_ (.A1(_0660_),
    .A2(_0665_),
    .B1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__a311o_1 _2309_ (.A1(_0660_),
    .A2(_0665_),
    .A3(_0666_),
    .B1(_0667_),
    .C1(_0661_),
    .X(_0668_));
 sky130_fd_sc_hd__xnor2_1 _2310_ (.A(_0663_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__a22o_1 _2311_ (.A1(_0624_),
    .A2(_0660_),
    .B1(_0637_),
    .B2(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__o21ba_1 _2312_ (.A1(_0637_),
    .A2(_0669_),
    .B1_N(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__xnor2_1 _2313_ (.A(_0657_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nor2_1 _2314_ (.A(_0608_),
    .B(_0672_),
    .Y(net22));
 sky130_fd_sc_hd__clkinv_2 _2315_ (.A(_0634_),
    .Y(_0673_));
 sky130_fd_sc_hd__mux2_1 _2316_ (.A0(_0607_),
    .A1(_0673_),
    .S(\A1.x[6] ),
    .X(_0674_));
 sky130_fd_sc_hd__a31o_1 _2317_ (.A1(_0611_),
    .A2(_0652_),
    .A3(_0637_),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__nand2_1 _2318_ (.A(_0660_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21a_1 _2319_ (.A1(_0607_),
    .A2(_0656_),
    .B1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _2320_ (.A(_0608_),
    .B(_0677_),
    .Y(net23));
 sky130_fd_sc_hd__and4b_1 _2321_ (.A_N(_0607_),
    .B(_0016_),
    .C(_0656_),
    .D(_0676_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _2322_ (.A(_0678_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _2323_ (.A(_0660_),
    .B(_0674_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _2324_ (.A(_0679_),
    .X(net16));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(\P1.qq[8] ),
    .A1(\P1.in[0] ),
    .S(net10),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _2326_ (.A(_0680_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _2327_ (.A(net15),
    .X(_0681_));
 sky130_fd_sc_hd__buf_4 _2328_ (.A(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__inv_2 _2329_ (.A(_0682_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _2330_ (.A(_0682_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _2331_ (.A(_0682_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _2332_ (.A(_0682_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _2333_ (.A(_0682_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _2334_ (.A(_0682_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _2335_ (.A(_0682_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _2336_ (.A(_0682_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _2337_ (.A(_0682_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _2338_ (.A(_0682_),
    .Y(_0026_));
 sky130_fd_sc_hd__buf_4 _2339_ (.A(_0681_),
    .X(_0683_));
 sky130_fd_sc_hd__inv_2 _2340_ (.A(_0683_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _2341_ (.A(_0683_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _2342_ (.A(_0683_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _2343_ (.A(_0683_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _2344_ (.A(_0683_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _2345_ (.A(_0683_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _2346_ (.A(_0683_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _2347_ (.A(_0683_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _2348_ (.A(_0683_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _2349_ (.A(_0683_),
    .Y(_0036_));
 sky130_fd_sc_hd__buf_4 _2350_ (.A(_0681_),
    .X(_0684_));
 sky130_fd_sc_hd__inv_2 _2351_ (.A(_0684_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _2352_ (.A(_0684_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _2353_ (.A(_0684_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _2354_ (.A(_0684_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _2355_ (.A(_0684_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _2356_ (.A(_0684_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _2357_ (.A(_0684_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _2358_ (.A(_0684_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _2359_ (.A(_0684_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _2360_ (.A(_0684_),
    .Y(_0046_));
 sky130_fd_sc_hd__buf_4 _2361_ (.A(_0681_),
    .X(_0685_));
 sky130_fd_sc_hd__inv_2 _2362_ (.A(_0685_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _2363_ (.A(_0685_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _2364_ (.A(_0685_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _2365_ (.A(_0685_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _2366_ (.A(_0685_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _2367_ (.A(_0685_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _2368_ (.A(_0685_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _2369_ (.A(_0685_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _2370_ (.A(_0685_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _2371_ (.A(_0685_),
    .Y(_0056_));
 sky130_fd_sc_hd__buf_4 _2372_ (.A(_0681_),
    .X(_0686_));
 sky130_fd_sc_hd__inv_2 _2373_ (.A(_0686_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _2374_ (.A(_0686_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _2375_ (.A(_0686_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _2376_ (.A(_0686_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _2377_ (.A(_0686_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _2378_ (.A(_0686_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _2379_ (.A(_0686_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _2380_ (.A(_0686_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _2381_ (.A(_0686_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _2382_ (.A(_0686_),
    .Y(_0066_));
 sky130_fd_sc_hd__buf_4 _2383_ (.A(_0629_),
    .X(_0687_));
 sky130_fd_sc_hd__inv_2 _2384_ (.A(_0687_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _2385_ (.A(_0687_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _2386_ (.A(_0687_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _2387_ (.A(_0687_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2388_ (.A(_0687_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _2389_ (.A(_0687_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _2390_ (.A(_0687_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _2391_ (.A(_0687_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _2392_ (.A(_0687_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _2393_ (.A(_0687_),
    .Y(_0076_));
 sky130_fd_sc_hd__buf_4 _2394_ (.A(_0629_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _2395_ (.A(_0688_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _2396_ (.A(_0688_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _2397_ (.A(_0688_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _2398_ (.A(_0688_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _2399_ (.A(_0688_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _2400_ (.A(_0688_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _2401_ (.A(_0688_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _2402_ (.A(_0688_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _2403_ (.A(_0688_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _2404_ (.A(_0688_),
    .Y(_0086_));
 sky130_fd_sc_hd__buf_4 _2405_ (.A(_0629_),
    .X(_0689_));
 sky130_fd_sc_hd__inv_2 _2406_ (.A(_0689_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _2407_ (.A(_0689_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2408_ (.A(_0689_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _2409_ (.A(_0689_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _2410_ (.A(_0689_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _2411_ (.A(_0689_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _2412_ (.A(_0689_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _2413_ (.A(_0689_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2414_ (.A(_0689_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _2415_ (.A(_0689_),
    .Y(_0096_));
 sky130_fd_sc_hd__buf_4 _2416_ (.A(_0629_),
    .X(_0690_));
 sky130_fd_sc_hd__inv_2 _2417_ (.A(_0690_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _2418_ (.A(_0690_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _2419_ (.A(_0690_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _2420_ (.A(_0690_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _2421_ (.A(_0690_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _2422_ (.A(_0690_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _2423_ (.A(_0690_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _2424_ (.A(_0690_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _2425_ (.A(_0690_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2426_ (.A(_0690_),
    .Y(_0106_));
 sky130_fd_sc_hd__buf_6 _2427_ (.A(_0629_),
    .X(_0691_));
 sky130_fd_sc_hd__inv_2 _2428_ (.A(_0691_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _2429_ (.A(_0691_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _2430_ (.A(_0691_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _2431_ (.A(_0691_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _2432_ (.A(_0691_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _2433_ (.A(_0691_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _2434_ (.A(_0691_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _2435_ (.A(_0691_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _2436_ (.A(_0691_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _2437_ (.A(_0691_),
    .Y(_0116_));
 sky130_fd_sc_hd__buf_4 _2438_ (.A(_0629_),
    .X(_0692_));
 sky130_fd_sc_hd__inv_2 _2439_ (.A(_0692_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _2440_ (.A(_0692_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _2441_ (.A(_0692_),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _2442_ (.A(_0692_),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _2443_ (.A(_0692_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _2444_ (.A(_0692_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _2445_ (.A(_0692_),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _2446_ (.A(_0692_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _2447_ (.A(_0692_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _2448_ (.A(_0692_),
    .Y(_0126_));
 sky130_fd_sc_hd__buf_6 _2449_ (.A(_0629_),
    .X(_0693_));
 sky130_fd_sc_hd__inv_2 _2450_ (.A(_0693_),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _2451_ (.A(_0693_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _2452_ (.A(_0693_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _2453_ (.A(_0693_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _2454_ (.A(_0693_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _2455_ (.A(_0693_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _2456_ (.A(_0693_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _2457_ (.A(_0693_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _2458_ (.A(_0693_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _2459_ (.A(_0693_),
    .Y(_0136_));
 sky130_fd_sc_hd__buf_4 _2460_ (.A(_0629_),
    .X(_0694_));
 sky130_fd_sc_hd__inv_2 _2461_ (.A(_0694_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(_0694_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _2463_ (.A(_0694_),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _2464_ (.A(_0694_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _2465_ (.A(_0694_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _2466_ (.A(_0694_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _2467_ (.A(_0694_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _2468_ (.A(_0694_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _2469_ (.A(_0694_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _2470_ (.A(_0694_),
    .Y(_0146_));
 sky130_fd_sc_hd__buf_4 _2471_ (.A(_0629_),
    .X(_0695_));
 sky130_fd_sc_hd__inv_2 _2472_ (.A(_0695_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _2473_ (.A(_0695_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _2474_ (.A(_0695_),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _2475_ (.A(_0695_),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _2476_ (.A(_0695_),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _2477_ (.A(_0695_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _2478_ (.A(_0695_),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _2479_ (.A(_0695_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _2480_ (.A(_0695_),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _2481_ (.A(_0695_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _2482_ (.A(_0681_),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _2483_ (.A(_0681_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _2484_ (.A(_0681_),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _2485_ (.A(_0681_),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _2486_ (.A(_0681_),
    .Y(_0161_));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(clknet_4_15_0_clk),
    .D(\m1.out[9] ),
    .Q(\P1.in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2488_ (.CLK(clknet_4_13_0_clk),
    .D(\m1.out[10] ),
    .Q(\P1.in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(clknet_4_15_0_clk),
    .D(\m1.out[11] ),
    .Q(\P1.in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(clknet_4_15_0_clk),
    .D(\m1.out[12] ),
    .Q(\P1.in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(clknet_4_12_0_clk),
    .D(\m1.out[13] ),
    .Q(\P1.in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(clknet_4_8_0_clk),
    .D(\m1.out[14] ),
    .Q(\P1.in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(clknet_4_8_0_clk),
    .D(\m1.out[15] ),
    .Q(\P1.in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(clknet_4_10_0_clk),
    .D(\m1.out[16] ),
    .Q(\P1.in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(clknet_4_9_0_clk),
    .D(\m2.out[9] ),
    .Q(\P1.in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(clknet_4_9_0_clk),
    .D(\m2.out[10] ),
    .Q(\P1.in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2497_ (.CLK(clknet_4_9_0_clk),
    .D(\m2.out[11] ),
    .Q(\P1.in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2498_ (.CLK(clknet_4_10_0_clk),
    .D(\m2.out[12] ),
    .Q(\P1.in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2499_ (.CLK(clknet_4_10_0_clk),
    .D(\m2.out[13] ),
    .Q(\P1.in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2500_ (.CLK(clknet_4_11_0_clk),
    .D(\m2.out[14] ),
    .Q(\P1.in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2501_ (.CLK(clknet_4_11_0_clk),
    .D(\m2.out[15] ),
    .Q(\P1.in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2502_ (.CLK(clknet_4_11_0_clk),
    .D(net48),
    .Q(\P1.in[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2503_ (.CLK(net11),
    .D(net2),
    .RESET_B(_0016_),
    .Q(\I1.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2504_ (.CLK(net11),
    .D(net3),
    .RESET_B(_0017_),
    .Q(\I1.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2505_ (.CLK(net11),
    .D(net4),
    .RESET_B(_0018_),
    .Q(\I1.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2506_ (.CLK(net11),
    .D(net5),
    .RESET_B(_0019_),
    .Q(\I1.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2507_ (.CLK(net11),
    .D(net6),
    .RESET_B(_0020_),
    .Q(\I1.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2508_ (.CLK(net11),
    .D(net7),
    .RESET_B(_0021_),
    .Q(\I1.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2509_ (.CLK(net11),
    .D(net8),
    .RESET_B(_0022_),
    .Q(\I1.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2510_ (.CLK(net11),
    .D(net9),
    .RESET_B(_0023_),
    .Q(\I1.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2511_ (.CLK(net12),
    .D(net2),
    .RESET_B(_0024_),
    .Q(\I2.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2512_ (.CLK(net12),
    .D(net3),
    .RESET_B(_0025_),
    .Q(\I2.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2513_ (.CLK(net12),
    .D(net4),
    .RESET_B(_0026_),
    .Q(\I2.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2514_ (.CLK(net12),
    .D(net5),
    .RESET_B(_0027_),
    .Q(\I2.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2515_ (.CLK(net12),
    .D(net6),
    .RESET_B(_0028_),
    .Q(\I2.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2516_ (.CLK(net12),
    .D(net7),
    .RESET_B(_0029_),
    .Q(\I2.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2517_ (.CLK(net12),
    .D(net8),
    .RESET_B(_0030_),
    .Q(\I2.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2518_ (.CLK(net12),
    .D(net9),
    .RESET_B(_0031_),
    .Q(\I2.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2519_ (.CLK(net13),
    .D(net2),
    .RESET_B(_0032_),
    .Q(\I3.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2520_ (.CLK(net13),
    .D(net3),
    .RESET_B(_0033_),
    .Q(\I3.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2521_ (.CLK(net13),
    .D(net4),
    .RESET_B(_0034_),
    .Q(\I3.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2522_ (.CLK(net13),
    .D(net5),
    .RESET_B(_0035_),
    .Q(\I3.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2523_ (.CLK(net13),
    .D(net6),
    .RESET_B(_0036_),
    .Q(\I3.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2524_ (.CLK(net13),
    .D(net7),
    .RESET_B(_0037_),
    .Q(\I3.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2525_ (.CLK(net13),
    .D(net8),
    .RESET_B(_0038_),
    .Q(\I3.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2526_ (.CLK(net13),
    .D(net9),
    .RESET_B(_0039_),
    .Q(\I3.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2527_ (.CLK(net14),
    .D(net2),
    .RESET_B(_0040_),
    .Q(\I4.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2528_ (.CLK(net14),
    .D(net3),
    .RESET_B(_0041_),
    .Q(\I4.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2529_ (.CLK(net14),
    .D(net4),
    .RESET_B(_0042_),
    .Q(\I4.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2530_ (.CLK(net14),
    .D(net5),
    .RESET_B(_0043_),
    .Q(\I4.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2531_ (.CLK(net14),
    .D(net6),
    .RESET_B(_0044_),
    .Q(\I4.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2532_ (.CLK(net14),
    .D(net7),
    .RESET_B(_0045_),
    .Q(\I4.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2533_ (.CLK(net14),
    .D(net8),
    .RESET_B(_0046_),
    .Q(\I4.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2534_ (.CLK(net14),
    .D(net9),
    .RESET_B(_0047_),
    .Q(\I4.out[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2535_ (.CLK(clknet_4_1_0_clk),
    .D(_0162_),
    .RESET_B(_0048_),
    .Q(\m1.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2536_ (.CLK(clknet_4_1_0_clk),
    .D(_0163_),
    .RESET_B(_0049_),
    .Q(\m1.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2537_ (.CLK(clknet_4_1_0_clk),
    .D(_0164_),
    .RESET_B(_0050_),
    .Q(\m1.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2538_ (.CLK(clknet_4_0_0_clk),
    .D(_0165_),
    .RESET_B(_0051_),
    .Q(\m1.b[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2539_ (.CLK(clknet_4_1_0_clk),
    .D(_0166_),
    .RESET_B(_0052_),
    .Q(\m1.b[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2540_ (.CLK(clknet_4_0_0_clk),
    .D(_0167_),
    .RESET_B(_0053_),
    .Q(\m1.b[5] ));
 sky130_fd_sc_hd__dfrtp_4 _2541_ (.CLK(clknet_4_0_0_clk),
    .D(_0168_),
    .RESET_B(_0054_),
    .Q(\m1.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2542_ (.CLK(clknet_4_0_0_clk),
    .D(_0169_),
    .RESET_B(_0055_),
    .Q(\m1.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2543_ (.CLK(clknet_4_3_0_clk),
    .D(_0170_),
    .RESET_B(_0056_),
    .Q(\m1.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2544_ (.CLK(clknet_4_4_0_clk),
    .D(_0171_),
    .RESET_B(_0057_),
    .Q(\m1.a[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2545_ (.CLK(clknet_4_1_0_clk),
    .D(_0172_),
    .RESET_B(_0058_),
    .Q(\m1.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2546_ (.CLK(clknet_4_4_0_clk),
    .D(_0173_),
    .RESET_B(_0059_),
    .Q(\m1.a[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2547_ (.CLK(clknet_4_4_0_clk),
    .D(_0174_),
    .RESET_B(_0060_),
    .Q(\m1.a[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2548_ (.CLK(clknet_4_0_0_clk),
    .D(_0175_),
    .RESET_B(_0061_),
    .Q(\m1.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2549_ (.CLK(clknet_4_0_0_clk),
    .D(_0176_),
    .RESET_B(_0062_),
    .Q(\m1.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2550_ (.CLK(clknet_4_1_0_clk),
    .D(_0177_),
    .RESET_B(_0063_),
    .Q(\m1.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2551_ (.CLK(clknet_4_3_0_clk),
    .D(_0178_),
    .RESET_B(_0064_),
    .Q(\m1.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2552_ (.CLK(clknet_4_6_0_clk),
    .D(_0179_),
    .RESET_B(_0065_),
    .Q(\m1.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2553_ (.CLK(clknet_4_5_0_clk),
    .D(_0180_),
    .RESET_B(_0066_),
    .Q(\m1.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2554_ (.CLK(clknet_4_7_0_clk),
    .D(_0181_),
    .RESET_B(_0067_),
    .Q(\m1.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2555_ (.CLK(clknet_4_7_0_clk),
    .D(_0182_),
    .RESET_B(_0068_),
    .Q(\m1.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2556_ (.CLK(clknet_4_13_0_clk),
    .D(_0183_),
    .RESET_B(_0069_),
    .Q(\m1.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2557_ (.CLK(clknet_4_7_0_clk),
    .D(_0184_),
    .RESET_B(_0070_),
    .Q(\m1.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2558_ (.CLK(clknet_4_7_0_clk),
    .D(_0185_),
    .RESET_B(_0071_),
    .Q(\m1.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2559_ (.CLK(clknet_4_7_0_clk),
    .D(_0186_),
    .RESET_B(_0072_),
    .Q(\m1.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2560_ (.CLK(clknet_4_15_0_clk),
    .D(_0187_),
    .RESET_B(_0073_),
    .Q(\m1.out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2561_ (.CLK(clknet_4_15_0_clk),
    .D(_0188_),
    .RESET_B(_0074_),
    .Q(\m1.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2562_ (.CLK(clknet_4_15_0_clk),
    .D(_0189_),
    .RESET_B(_0075_),
    .Q(\m1.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2563_ (.CLK(clknet_4_15_0_clk),
    .D(_0190_),
    .RESET_B(_0076_),
    .Q(\m1.out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2564_ (.CLK(clknet_4_12_0_clk),
    .D(_0191_),
    .RESET_B(_0077_),
    .Q(\m1.out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2565_ (.CLK(clknet_4_12_0_clk),
    .D(_0192_),
    .RESET_B(_0078_),
    .Q(\m1.out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2566_ (.CLK(clknet_4_6_0_clk),
    .D(_0193_),
    .RESET_B(_0079_),
    .Q(\m1.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2567_ (.CLK(clknet_4_12_0_clk),
    .D(_0194_),
    .RESET_B(_0080_),
    .Q(\m1.out[16] ));
 sky130_fd_sc_hd__dfrtp_2 _2568_ (.CLK(clknet_4_2_0_clk),
    .D(_0195_),
    .RESET_B(_0081_),
    .Q(\m2.b[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2569_ (.CLK(clknet_4_2_0_clk),
    .D(_0196_),
    .RESET_B(_0082_),
    .Q(\m2.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2570_ (.CLK(clknet_4_2_0_clk),
    .D(_0197_),
    .RESET_B(_0083_),
    .Q(\m2.b[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2571_ (.CLK(clknet_4_3_0_clk),
    .D(_0198_),
    .RESET_B(_0084_),
    .Q(\m2.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2572_ (.CLK(clknet_4_2_0_clk),
    .D(_0199_),
    .RESET_B(_0085_),
    .Q(\m2.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2573_ (.CLK(clknet_4_2_0_clk),
    .D(_0200_),
    .RESET_B(_0086_),
    .Q(\m2.b[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2574_ (.CLK(clknet_4_2_0_clk),
    .D(_0201_),
    .RESET_B(_0087_),
    .Q(\m2.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2575_ (.CLK(clknet_4_2_0_clk),
    .D(_0202_),
    .RESET_B(_0088_),
    .Q(\m2.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2576_ (.CLK(clknet_4_3_0_clk),
    .D(_0203_),
    .RESET_B(_0089_),
    .Q(\m2.a[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2577_ (.CLK(clknet_4_3_0_clk),
    .D(_0204_),
    .RESET_B(_0090_),
    .Q(\m2.a[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2578_ (.CLK(clknet_4_3_0_clk),
    .D(_0205_),
    .RESET_B(_0091_),
    .Q(\m2.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2579_ (.CLK(clknet_4_2_0_clk),
    .D(_0206_),
    .RESET_B(_0092_),
    .Q(\m2.a[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2580_ (.CLK(clknet_4_2_0_clk),
    .D(_0207_),
    .RESET_B(_0093_),
    .Q(\m2.a[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2581_ (.CLK(clknet_4_2_0_clk),
    .D(_0208_),
    .RESET_B(_0094_),
    .Q(\m2.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2582_ (.CLK(clknet_4_2_0_clk),
    .D(_0209_),
    .RESET_B(_0095_),
    .Q(\m2.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2583_ (.CLK(clknet_4_2_0_clk),
    .D(_0210_),
    .RESET_B(_0096_),
    .Q(\m2.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2584_ (.CLK(clknet_4_14_0_clk),
    .D(_0211_),
    .RESET_B(_0097_),
    .Q(\m2.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2585_ (.CLK(clknet_4_13_0_clk),
    .D(_0212_),
    .RESET_B(_0098_),
    .Q(\m2.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2586_ (.CLK(clknet_4_13_0_clk),
    .D(_0213_),
    .RESET_B(_0099_),
    .Q(\m2.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2587_ (.CLK(clknet_4_13_0_clk),
    .D(_0214_),
    .RESET_B(_0100_),
    .Q(\m2.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2588_ (.CLK(clknet_4_15_0_clk),
    .D(_0215_),
    .RESET_B(_0101_),
    .Q(\m2.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2589_ (.CLK(clknet_4_14_0_clk),
    .D(_0216_),
    .RESET_B(_0102_),
    .Q(\m2.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2590_ (.CLK(clknet_4_14_0_clk),
    .D(_0217_),
    .RESET_B(_0103_),
    .Q(\m2.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2591_ (.CLK(clknet_4_8_0_clk),
    .D(_0218_),
    .RESET_B(_0104_),
    .Q(\m2.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2592_ (.CLK(clknet_4_8_0_clk),
    .D(_0219_),
    .RESET_B(_0105_),
    .Q(\m2.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2593_ (.CLK(clknet_4_8_0_clk),
    .D(_0220_),
    .RESET_B(_0106_),
    .Q(\m2.out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2594_ (.CLK(clknet_4_9_0_clk),
    .D(_0221_),
    .RESET_B(_0107_),
    .Q(\m2.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2595_ (.CLK(clknet_4_9_0_clk),
    .D(_0222_),
    .RESET_B(_0108_),
    .Q(\m2.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2596_ (.CLK(clknet_4_10_0_clk),
    .D(_0223_),
    .RESET_B(_0109_),
    .Q(\m2.out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2597_ (.CLK(clknet_4_10_0_clk),
    .D(_0224_),
    .RESET_B(_0110_),
    .Q(\m2.out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2598_ (.CLK(clknet_4_11_0_clk),
    .D(_0225_),
    .RESET_B(_0111_),
    .Q(\m2.out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2599_ (.CLK(clknet_4_11_0_clk),
    .D(_0226_),
    .RESET_B(_0112_),
    .Q(\m2.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2600_ (.CLK(clknet_4_10_0_clk),
    .D(_0227_),
    .RESET_B(_0113_),
    .Q(\m2.out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2601_ (.CLK(clknet_4_6_0_clk),
    .D(_0228_),
    .RESET_B(_0114_),
    .Q(\m1.multa_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2602_ (.CLK(clknet_4_6_0_clk),
    .D(_0229_),
    .RESET_B(_0115_),
    .Q(\m1.multa_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2603_ (.CLK(clknet_4_4_0_clk),
    .D(_0230_),
    .RESET_B(_0116_),
    .Q(\m1.multa_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2604_ (.CLK(clknet_4_6_0_clk),
    .D(_0231_),
    .RESET_B(_0117_),
    .Q(\m1.multa_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2605_ (.CLK(clknet_4_7_0_clk),
    .D(_0232_),
    .RESET_B(_0118_),
    .Q(\m1.multa_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2606_ (.CLK(clknet_4_7_0_clk),
    .D(_0233_),
    .RESET_B(_0119_),
    .Q(\m1.multa_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2607_ (.CLK(clknet_4_7_0_clk),
    .D(_0234_),
    .RESET_B(_0120_),
    .Q(\m1.multa_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2608_ (.CLK(clknet_4_7_0_clk),
    .D(_0235_),
    .RESET_B(_0121_),
    .Q(\m1.multa_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2609_ (.CLK(clknet_4_5_0_clk),
    .D(_0236_),
    .RESET_B(_0122_),
    .Q(\m1.multa_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2610_ (.CLK(clknet_4_5_0_clk),
    .D(_0237_),
    .RESET_B(_0123_),
    .Q(\m1.multa_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2611_ (.CLK(clknet_4_5_0_clk),
    .D(_0238_),
    .RESET_B(_0124_),
    .Q(\m1.multa_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2612_ (.CLK(clknet_4_5_0_clk),
    .D(_0239_),
    .RESET_B(_0125_),
    .Q(\m1.multa_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2613_ (.CLK(clknet_4_5_0_clk),
    .D(_0240_),
    .RESET_B(_0126_),
    .Q(\m1.multa_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2614_ (.CLK(clknet_4_6_0_clk),
    .D(_0241_),
    .RESET_B(_0127_),
    .Q(\m1.multa_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2615_ (.CLK(clknet_4_3_0_clk),
    .D(_0242_),
    .RESET_B(_0128_),
    .Q(\m1.multa_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2616_ (.CLK(clknet_4_0_0_clk),
    .D(_0243_),
    .RESET_B(_0129_),
    .Q(\m1.multa_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2617_ (.CLK(clknet_4_10_0_clk),
    .D(_0000_),
    .RESET_B(_0130_),
    .Q(\A1.x[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2618_ (.CLK(clknet_4_11_0_clk),
    .D(_0007_),
    .RESET_B(_0131_),
    .Q(\A1.x[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2619_ (.CLK(clknet_4_10_0_clk),
    .D(_0008_),
    .RESET_B(_0132_),
    .Q(\A1.x[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2620_ (.CLK(clknet_4_11_0_clk),
    .D(_0009_),
    .RESET_B(_0133_),
    .Q(\A1.x[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2621_ (.CLK(clknet_4_11_0_clk),
    .D(_0010_),
    .RESET_B(_0134_),
    .Q(\A1.x[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2622_ (.CLK(clknet_4_11_0_clk),
    .D(_0011_),
    .RESET_B(_0135_),
    .Q(\A1.x[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2623_ (.CLK(clknet_4_11_0_clk),
    .D(_0012_),
    .RESET_B(_0136_),
    .Q(\A1.x[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2624_ (.CLK(clknet_4_11_0_clk),
    .D(_0013_),
    .RESET_B(_0137_),
    .Q(\A1.x[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2625_ (.CLK(clknet_4_8_0_clk),
    .D(_0014_),
    .RESET_B(_0138_),
    .Q(\P1.qq[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2626_ (.CLK(clknet_4_9_0_clk),
    .D(_0015_),
    .RESET_B(_0139_),
    .Q(\P1.qq[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2627_ (.CLK(clknet_4_9_0_clk),
    .D(_0001_),
    .RESET_B(_0140_),
    .Q(\P1.qq[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2628_ (.CLK(clknet_4_9_0_clk),
    .D(_0002_),
    .RESET_B(_0141_),
    .Q(\P1.qq[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2629_ (.CLK(clknet_4_9_0_clk),
    .D(_0003_),
    .RESET_B(_0142_),
    .Q(\P1.qq[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2630_ (.CLK(clknet_4_9_0_clk),
    .D(_0004_),
    .RESET_B(_0143_),
    .Q(\P1.qq[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2631_ (.CLK(clknet_4_10_0_clk),
    .D(_0005_),
    .RESET_B(_0144_),
    .Q(\P1.qq[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2632_ (.CLK(clknet_4_8_0_clk),
    .D(_0006_),
    .RESET_B(_0145_),
    .Q(\P1.qq[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2633_ (.CLK(clknet_4_12_0_clk),
    .D(_0244_),
    .RESET_B(_0146_),
    .Q(\m2.multa_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2634_ (.CLK(clknet_4_13_0_clk),
    .D(_0245_),
    .RESET_B(_0147_),
    .Q(\m2.multa_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2635_ (.CLK(clknet_4_12_0_clk),
    .D(_0246_),
    .RESET_B(_0148_),
    .Q(\m2.multa_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2636_ (.CLK(clknet_4_15_0_clk),
    .D(_0247_),
    .RESET_B(_0149_),
    .Q(\m2.multa_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2637_ (.CLK(clknet_4_13_0_clk),
    .D(_0248_),
    .RESET_B(_0150_),
    .Q(\m2.multa_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2638_ (.CLK(clknet_4_14_0_clk),
    .D(_0249_),
    .RESET_B(_0151_),
    .Q(\m2.multa_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2639_ (.CLK(clknet_4_14_0_clk),
    .D(_0250_),
    .RESET_B(_0152_),
    .Q(\m2.multa_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2640_ (.CLK(clknet_4_14_0_clk),
    .D(_0251_),
    .RESET_B(_0153_),
    .Q(\m2.multa_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2641_ (.CLK(clknet_4_14_0_clk),
    .D(_0252_),
    .RESET_B(_0154_),
    .Q(\m2.multa_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2642_ (.CLK(clknet_4_14_0_clk),
    .D(_0253_),
    .RESET_B(_0155_),
    .Q(\m2.multa_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2643_ (.CLK(clknet_4_8_0_clk),
    .D(_0254_),
    .RESET_B(_0156_),
    .Q(\m2.multa_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2644_ (.CLK(clknet_4_10_0_clk),
    .D(_0255_),
    .RESET_B(_0157_),
    .Q(\m2.multa_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2645_ (.CLK(clknet_4_11_0_clk),
    .D(_0256_),
    .RESET_B(_0158_),
    .Q(\m2.multa_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2646_ (.CLK(clknet_4_11_0_clk),
    .D(_0257_),
    .RESET_B(_0159_),
    .Q(\m2.multa_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2647_ (.CLK(clknet_4_11_0_clk),
    .D(_0258_),
    .RESET_B(_0160_),
    .Q(\m2.multa_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2648_ (.CLK(clknet_4_11_0_clk),
    .D(_0259_),
    .RESET_B(_0161_),
    .Q(\m2.multa_reg[15] ));
 sky130_fd_sc_hd__conb_1 mac_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 mac_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 mac_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 mac_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 mac_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 mac_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 mac_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 mac_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 mac_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 mac_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 mac_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 mac_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 mac_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 mac_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 mac_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 mac_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 mac_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 mac_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 mac_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 mac_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 mac_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 mac_47 (.LO(net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(clken),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(in[4]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(in[5]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(ld),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(ld1),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(ld2),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(ld3),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(ld4),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(rst),
    .X(net15));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(out[10]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(out[5]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(out[7]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(out[8]));
 sky130_fd_sc_hd__conb_1 mac_25 (.LO(net25));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\m2.out[16] ),
    .X(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__B (.DIODE(\P1.in[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__RESET_B (.DIODE(_0016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__B (.DIODE(_0016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__B2 (.DIODE(_0016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B (.DIODE(_0016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__B (.DIODE(_0330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__S (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__S (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__S (.DIODE(_0544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__S (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__B (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A0 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__B2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__B2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A0 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__B2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__A0 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__A2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__A2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__C (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__A0 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__A2 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__A0 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__B2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__A0 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__C (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__C (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__B1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__D (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A0 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__B2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A0 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__B2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__A1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__A1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__A0 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A2_N (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__D (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1366__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__A2 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__C (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A0 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A2 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__C (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A2 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__C (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A2 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__B1 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1334__C (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__B (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__D (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A0 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__B2 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A1 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__A1 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__A1 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A0 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__C (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__D (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__B1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__D (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__D (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__B1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1334__D (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__A0 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B2 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__B2 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__B (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__A0 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A1_N (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__B (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__B1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__C1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__S (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__C1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__B1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__B (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__B (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__B (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1554__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__C (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__S (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__S (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A0 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__C (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__D (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A0 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__C (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__C (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A2 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__B1 (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__B (.DIODE(_1038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A0 (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__B (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__B (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__B1 (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__D (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__B1 (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__B (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__B1 (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A2 (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__B (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__A0 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A2 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__C (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__A2 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A2 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A2 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__B1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__C (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__B (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__D (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__A0 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__B2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__B2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__B (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__A (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__A1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__A (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__A1 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__B (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A1 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__B (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__A (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A0 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__A (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A0 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__B2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__A (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__A (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__B2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__B (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__A (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A1 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A0 (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__B (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A1 (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__A (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A1_N (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__B (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A1 (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__B1 (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__A (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(clken));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(ld));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(ld1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(ld2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(ld3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(ld4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A2 (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__C1 (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__B (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__B (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__A (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__A (.DIODE(\m1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__D (.DIODE(\m1.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__A0 (.DIODE(\m1.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__B (.DIODE(\m1.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__B (.DIODE(\m1.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__D (.DIODE(\m1.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__A0 (.DIODE(\m1.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__B (.DIODE(\m1.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__B (.DIODE(\m1.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__S (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__CLK (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__CLK (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1928 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1917 ();
 assign io_oeb[0] = net25;
 assign io_oeb[10] = net35;
 assign io_oeb[11] = net36;
 assign io_oeb[12] = net37;
 assign io_oeb[13] = net38;
 assign io_oeb[14] = net39;
 assign io_oeb[15] = net40;
 assign io_oeb[1] = net26;
 assign io_oeb[2] = net27;
 assign io_oeb[3] = net28;
 assign io_oeb[4] = net29;
 assign io_oeb[5] = net30;
 assign io_oeb[6] = net31;
 assign io_oeb[7] = net32;
 assign io_oeb[8] = net33;
 assign io_oeb[9] = net34;
 assign out[0] = net41;
 assign out[11] = net46;
 assign out[12] = net45;
 assign out[13] = net44;
 assign out[14] = net43;
 assign out[15] = net42;
 assign out[9] = net47;
endmodule

