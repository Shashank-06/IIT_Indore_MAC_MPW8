magic
tech sky130A
magscale 1 2
timestamp 1671540496
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1436 178848 117552
<< metal2 >>
rect 3422 0 3478 800
rect 7102 0 7158 800
rect 10782 0 10838 800
rect 14462 0 14518 800
rect 18142 0 18198 800
rect 21822 0 21878 800
rect 25502 0 25558 800
rect 29182 0 29238 800
rect 32862 0 32918 800
rect 36542 0 36598 800
rect 40222 0 40278 800
rect 43902 0 43958 800
rect 47582 0 47638 800
rect 51262 0 51318 800
rect 54942 0 54998 800
rect 58622 0 58678 800
rect 62302 0 62358 800
rect 65982 0 66038 800
rect 69662 0 69718 800
rect 73342 0 73398 800
rect 77022 0 77078 800
rect 80702 0 80758 800
rect 84382 0 84438 800
rect 88062 0 88118 800
rect 91742 0 91798 800
rect 95422 0 95478 800
rect 99102 0 99158 800
rect 102782 0 102838 800
rect 106462 0 106518 800
rect 110142 0 110198 800
rect 113822 0 113878 800
rect 117502 0 117558 800
rect 121182 0 121238 800
rect 124862 0 124918 800
rect 128542 0 128598 800
rect 132222 0 132278 800
rect 135902 0 135958 800
rect 139582 0 139638 800
rect 143262 0 143318 800
rect 146942 0 146998 800
rect 150622 0 150678 800
rect 154302 0 154358 800
rect 157982 0 158038 800
rect 161662 0 161718 800
rect 165342 0 165398 800
rect 169022 0 169078 800
rect 172702 0 172758 800
rect 176382 0 176438 800
<< obsm2 >>
rect 3424 856 176436 117541
rect 3534 800 7046 856
rect 7214 800 10726 856
rect 10894 800 14406 856
rect 14574 800 18086 856
rect 18254 800 21766 856
rect 21934 800 25446 856
rect 25614 800 29126 856
rect 29294 800 32806 856
rect 32974 800 36486 856
rect 36654 800 40166 856
rect 40334 800 43846 856
rect 44014 800 47526 856
rect 47694 800 51206 856
rect 51374 800 54886 856
rect 55054 800 58566 856
rect 58734 800 62246 856
rect 62414 800 65926 856
rect 66094 800 69606 856
rect 69774 800 73286 856
rect 73454 800 76966 856
rect 77134 800 80646 856
rect 80814 800 84326 856
rect 84494 800 88006 856
rect 88174 800 91686 856
rect 91854 800 95366 856
rect 95534 800 99046 856
rect 99214 800 102726 856
rect 102894 800 106406 856
rect 106574 800 110086 856
rect 110254 800 113766 856
rect 113934 800 117446 856
rect 117614 800 121126 856
rect 121294 800 124806 856
rect 124974 800 128486 856
rect 128654 800 132166 856
rect 132334 800 135846 856
rect 136014 800 139526 856
rect 139694 800 143206 856
rect 143374 800 146886 856
rect 147054 800 150566 856
rect 150734 800 154246 856
rect 154414 800 157926 856
rect 158094 800 161606 856
rect 161774 800 165286 856
rect 165454 800 168966 856
rect 169134 800 172646 856
rect 172814 800 176326 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 32862 0 32918 800 6 clk
port 1 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 clken
port 2 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 in[0]
port 3 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 in[1]
port 4 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 in[2]
port 5 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 in[3]
port 6 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 in[4]
port 7 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 in[5]
port 8 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 in[6]
port 9 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 in[7]
port 10 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 io_oeb[0]
port 11 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 io_oeb[10]
port 12 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 io_oeb[11]
port 13 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 io_oeb[12]
port 14 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 io_oeb[13]
port 15 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 io_oeb[14]
port 16 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 io_oeb[15]
port 17 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 io_oeb[1]
port 18 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 io_oeb[2]
port 19 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 io_oeb[3]
port 20 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 io_oeb[4]
port 21 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 io_oeb[5]
port 22 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 io_oeb[6]
port 23 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 io_oeb[7]
port 24 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 io_oeb[8]
port 25 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 io_oeb[9]
port 26 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 ld
port 27 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 ld1
port 28 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 ld2
port 29 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 ld3
port 30 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 ld4
port 31 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 out[0]
port 32 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 out[10]
port 33 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 out[11]
port 34 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 out[12]
port 35 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 out[13]
port 36 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 out[14]
port 37 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 out[15]
port 38 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 out[1]
port 39 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 out[2]
port 40 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 out[3]
port 41 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 out[4]
port 42 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 out[5]
port 43 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 out[6]
port 44 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 out[7]
port 45 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 out[8]
port 46 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 out[9]
port 47 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 rst
port 48 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 50 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9340936
string GDS_FILE /home/sky/MPW8/IIT_Indore_MAC_MPW8/openlane/mac/runs/22_12_20_04_43/results/signoff/mac.magic.gds
string GDS_START 493950
<< end >>

